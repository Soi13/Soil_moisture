PK   �p1Y��O�K  ��     cirkitFile.json�]�o�8�W�W�Ib{��a�
�=$�!Kr�[���r�{E��#)َ,Qg&m�pyhq8�8����Y�~*��lW�OE�/w��S��CZ���W����.���c�>=�n�ؿ��ϧ"�v�O�m���L��Vk���4X�qZdL1V�/����P�TgR��:(�PRI�i�
2�E����+�djv?������q����uW���{���k�"�pp�g�C�:kԼ�{�!7�uK�fL��8r�2�Fe�g�t��Y΋��<	�J�A�,�2��U�y���+r�3�6g��!�?ֿp���Y���Fy �(
t�V�*�<�V\$����㶛D�-Qc��
56G������8r�q�v�������@������ ��!4�߽���1�cu�	j��B` 6<44��l_�	�0��7rw3�+�z��>_
����}��0c�|)0-�������}��-v��Ԡ�{xl��{oPw��u�{o�E8���?�g��2 �;bpH��C��: c�m��S������)s��6�
����5,d��� ��5Z�B'�"H�H-�DKD�%&ђ�hэ��Ġ΁w��".0jh��h��~5��l�QC`F�`� �	�2�33M�z!�"nQ�+�QӲpZ��&w(�x��5FM��d�1��4D�iP�iP�'QM�h��04H�e2��&��
��Z&Y��#��Ы�i.=;���r�,�x  N�Lf:� ����
���Np�i���y��s8'48��;��14�2h�@�$uBS1�M��EME��D��\��-�6fO�i�	!��zs�s�:�lnc[�*� sx-�D� �"I�(-���DKB�EӠ��4�e4�e4�e4 f4f4f4f4 f4(�4(�DL�bN�bN�bN�bN�bN�bN�b>�bpn�e���^�$�����I��sx-���6�Zh�;G�sjh�;G�sjh<G�sj&A�m�L����k��8���2	<pn�e�F��^˴������6�:7��Q7U�2�cvâ��sY���&͊|Yn��*/���-�*���9�>c8�Ш����5��V���,�3fh�b>E��D}z���L�\�+/K���r���3��X�;��
��PG��J�t���q�耾W���4��ơ^ s:GfhC��Ǡ�*w�LԘn� ��L�w��~Q%~��?l�I��Pst�$��� x�g��?	��C�P�F��6p`�f@��&hi�;�`�1|���h�@��,����G�5@�F�vD��0���j/`��S��"	��=L�Z�F/��%%aO�S@4	4��iO�i���.���n��ۢ�C�cK6��ǭ�k7�ȪML��/�����#�'���'乭�scX|2,@]%����y,b�����P���b�aA�j1Q,b�y����y� �-�(�j1/�a>��2/��rVX"�Xs,����U���#W^b����jˋ���Fx\p���w&�������B���ë0	�78�1a�Ȅ(�4�B� 7@Ȟ��X�B��l`;� ��:N�����#���쮆�<�囘�����1�@k71�Ǭ�׼X�/ nb�3`fk7�j���:���Mv@���/kb�Z�df	Ғ���<����ɬ$��.�Ŭ0��.��?��.���w�m�~u	P����=���ݻ!4�J�6�Cv�t� `�ƚ�ƈۢ�6\6�t���/��}��{+%�=�Je���nO������MT`�r�no�ń�BɾGĽW;ُ>q/�E�S��k����������Ȣ�~�z5(��h�^L�z~v�s����&]��.��p��_��h�ڦ���Mq�)i��~k�X�)l��~�h�D�I�M�ߤ�&�o�m��5��4�/f���f���4_��ʖW�w�M������r2����N͵/���j�TTuY��Ѿ�d�/k�}\�"���j.$_�R��h����I%��E�"F�u bY�q��
�:Ց��i��N_ 6��X�N�Y���g��4Z�fz�Ó�]V٦h�薫x�撅��[��Z��x!��ED�*��.�+��$::]NM��i����x!��B(N}b'���-��D�U���A�n\��G�7�!kE�c���qǗ�J*�N�%#7~���ڟc_�>�~!�X��X-dl.�V8n��ʅ��K��8��v�C���G�5
��� N�i�DFǋ��Qd@�\��݄"��}wf,���xP�֌kP��Ϛ��G̴�]�y)~�O�x�ݧJ��-6�ąfzd!������?ԇ�ܝ6�-�B ������g��H���~4[t�>ڿm�|�)��_o޽	��.�tؖ��f������ߌ���:��Ӹ/���}���kU�CY�9��P�zL��u�Շ��Ʀ�\�<�Oi���[��t	Ԯ�[R�n�x��Z4;�]��|�X,t�� gl(�� a!���T�Rz�RM�)�0�S�3�O#�H��=l������æ%:_�{7{l�Za�S#�B?�9���ϳKL������$�m��z���:79�>t�bC�? 6�b��h��@��������y��Ͽ��0�?�ƗD�d��'n���;^��]q,��f2`y�+��`�M�]�����#���	P��6ޙ3e&y����0���`�R|�̸E�ƍj�,�[���7#��"�XʊER%��$f��z�c�t���\
�x���7�,$�
����[�>��!Ɗ�7'~�Z�-J{��Z|���iy��6w��wO�%l�P�kk_����?�y�`OkG�7���フ���
�c��~v4��i�P�oN'��UQ��V��a?�g�
_�f�ew�����u�f�;Դ�ߗ۷�kzq�)+���*`J����(�f��L8��]��ߧ��S����nf�����m������ͭ������Ҝ���B+0�:��n0 u��n�� �k��5ƔFg�V���Έ������#f����@�sp���ѓ�o�����_])����L�tj�HOH�y�:%�4!�D� Ҵ��@ݜ�@"Q n��:L�`�����04�ߓr� �FBM.�ɋ��{c�)�|럥XB0)�t!e�B���BhPJ1�q*0�x8¹pP=)]��$�����$	�^�AS��J@R��WOH�b�����9��bri���ӻ6v9=�s�q~��1煔�j��k�B��:��h����D0`�����N|z��I:�}������������+R���F$5aG#�E�qz�?�R�p��t2)0����M�ɕR���]���UOj��w���Q�QP�Q��Q������,���C�Pݬ/L*&����J��So1
Ǟ���7��QS�Q��4�誙F�x)5�BJt�0�(m���R�\�1���Iñ��: a��th���S���y�O]��<?|��Bj����$�K]�	)�c�ݔP��j���sE�w�Ԩ��(��+� υ�0�(�� B>G�'�e[ Pn6�ֿ�uQ��f?��xڻ?��/���n������������S��g��?��*��҈��� PK   �p1Y8�w���  ��  /   images/0392a38f-5b07-422b-a303-6a624800f9c8.pngt�eT]ݒ6�qww���=����7���N$xpw���!���s�����������%O�ڟ�eP	A ����*�A���#���'@��,��)F��A\R&�	ܥ��՜,ݽL\-@^^^,6�vnf&�,N�V'�� 9HNRL�;�軗7��@G��#WX���&$2RU=
�(�h�OLR���
	B�X�*�>�z�hP��2���H���;�G/��Ga�������0UD#�� �|y)_k%�E�	n!|�Q�xH��:o�'
�󊳡k���AV��Ehl�atܽ�V�}�-£�z��4*�����R��[C��sN,�4����t�P��P1�s��k�a��[��9Uӳ��$ceoZ���Hd��nD�N���z]`bX��;��n>��v���*/2��Ю+D�Ѕf2g��
ZU#��*�*�Ɏ�$�r\�gq+�R]�P��blz��r"�V�m�BO���N�J�Ӕ1>��Ptǟ��.�;���r84(#!*&S�����C�,�g�"��oá�l�mI�b��k�}�*[�:���rF�չ&�!O1ogX���@*�n��^i���KtW�U�,�p��d��v+�)tpʊ��мb�!�2�L��uh<�V?y�M P��<�	���?Sby�J������Hb��<խ:9�c��Qv|З�͉�c
�:���9�	�(���)HBOT�����p-��b��A�Aa���b��HȣqH�_�ۃ�#J��s�'��L�	B�r6���ul4{��x��i����=8�O�\QF	A�|�&�
>�9�Kv�mb�U��tbDev;ORq�`�o�Y����v�G�P��ˡ���h�3irq2��[�&�����l ��E�lP�骟Mߑ�J��2��E���b�RE��/��m�*�t�jz�Ƞ�*�M�'.a�+F0�6@��.g,S�P�xZ ^rߍ�!*���,�)e�q}	�z�"y�L�bTtE�Bs��$g.������u⾂)c���.ȉ@�F���t�>�b�XC��433�024rQ�I��ʑ��������H���L8�X�o\�8�qgt�w�t��|h7��*�� 	�O���bcP�����?y$S�>���Gb�gT2R��dܕ�u��|F�S`��Gz��)K�jY^��2��Fl������\���o\��8�\G�!�1&h�A�����m�"5��#��
�A��x���+n�<X~&Aڷ�cQ���V!'�졅��rx��}�Elv�4{↽) ����o+~i��K�#\�o�XF#��`�kL����0�TO-�;����"�Ck�������G�f����`b/ ��M��vgC�1|���Ou+�����ܕ�+nR�Q�1�.��7 f ��̫Č_��zE�E7�bc��v�ɑ�*�j	n�g�_&8s�S�J\Y`4`��J����g5%e����5�
D�6'9�eS!�G0���s��s�~�ԗd*@���%	� �[��J���0��)�nV���ݪ4UY$���G��6)���Tư�:�&�X?Ƌ�j����^�bs�7ߺ
J�M�i�S�ZV�:h�+zO�8�֕e�8DlF0�}G�SM.=4)r�1Mw�7��S2��Hb��)UG��>b#
��+0�B��6ϸ�������Y���Q�I��F�b�O��&�Y#
忶�&�A4Պ�@퉲��%�̇���5(b���(����7_�,�r��w[|�6�.$��W["3-��������'27DMbɥGg"yS�&�A(�3`qe�Qѩ�,?��ol
�Mb�KN�P�B��L�V���]Y �@�q"׬���p� �Lg�6gn�::$���/n�(��SʒĴ42��FE}VXD) QJ�|� �7�J&tQ��F>m�wzȥgg"��$�C�5	�:4iF��6/�$r��H{��3p�H�M���T���n^���ռ3 ��'C�h��GT�`�i��m�C
F7�;�V�~_f���BV�?�䪜B9����[�Ҝ������B�t���a܅�oV�ҷqi�t���a؅�%۬��/Z�-����:�B��/�֨�`q�{`9���@��"�k꿚��]�w�����C��0����$F��}�I����·�T��Qs�6M�C1��sX�n��V ��M��Bz�5���&�"\�/}Oto��#�ŋo�x4�3SHI��oWC=�/��@p�r�5�4�{f:�Yᖧ�d"�r4+���({I� | �B �!�{8��;�>��X�@;��Z,��l�qp�.����+����VR&���T�vL�Ц�ۅ���N�<��ٗOt^|g@������s�<�
�K�\�*���VT&�̿��,�F�ㆹ�-�P��4���:��Hy��e�=��f��Y���Vκ�f[j�!�Y<�&�}�R��u�r������V�v�Rݩ�����Ue�Yeu �d�R�{g`���y.�ddd��H��=�s����=q8���^�"l,��R���FJ�@?m��a\��-a*��T*ӛոe�:���:�
p�Z��A�f��T�]Hj�b���T@��1 �ah�i�d"�������3��h����_�|x���o��D�_�Ə��*>KR��뱖CJ�$2��v��fX�4�S}�Q:Q��:pEsR�#c\M�5�2k�̰�CK���������m|+'�dQ���^�(�r";E����;:���E�8j{�4Qsz $M�G�j�@�ä9�ˬ�Y	�׵�w��z�׾���>��h���;�Y'�(ݕ�Q�1gJ���,7f�O��g<C.��$d�� OǋG������Rl���f\m)ts�F��O���s��֥8=�҆�w6 ���]s�6���>�<|h�^��>�R�7.`(��a���gf\�����Rl"�V�D�J��Qh�1�<��֊̰Je��8��1�f��<�mUEH�'W�]er�X�A��hv���N��B9��vWC��i���N�12�X*�f�J���.�����ԩ+��N�cN+��KG#î�t���%��5T�����?�t�$CW�n	(��-�z�L�OѼ.��ƕ1�������(�Q^(}��v��I���(/�-c- 9�?y�]��ha?�R���+3����'�>ﰸ���d���z�a����^=�,�k� AP �W,��:O�7dcrP��8.^j�9>2lh�1�/	x����V
ퟛM�J�����.}񈌓�A"� �0Ɂ�^��U�3z���s������
�7���L������.CF���*�Ġ�Vc�儬vݔsZ��R$�2����`��3� g�)��� 敜�[�����^�3�<AL�J��r�ވG�G�>Ձ�ߴ���l)O�mJҷ,��v� >�z.Fe[$o�s<�F�,�xL��̾����}}��6�q	5����%��1��ŵ�4���=�HB��^%�m�������ԫ��~��ch5�՛�%��YCY펈��X���]�łM�&�"$�,��?�E��.����)��V���4R�\�nӱ�N���l��Nz�h77DȚ�����>9ѫ��߹���F��|�Q���ex!��z*�=
$��_� �y�tʹ�ǈ�Q�L	y�T�sNi�9��Ґ� �yM�7��)O;���)�̲�߽(&'�������W��;f�����=�`A�ivj�=KAͻ5����t���-P�G�:d�f`,��y��Wߞ�U l�x�;Eؗ��`c��(�q�ÕL������Cp5�7��q�E���4�e��F�R��P7�ݚ!U�h�Zz�c�����\���c��?v�cm|��������b^�_�zG��_���5泩�][5��q�J�.VVˣ��A��Q�~F���5��������+�,y/�N;�C1�XSLf/&�&�}��E���V��`��ow6wn��vj��ߚ̳ 8���[O���lԼ_F�%m�[y�U\��K/�u��FXAξ�S�^��xA��F��;��Ki�M�[U��۸#��j�$�mE=ul���Ҏjg�2hɶ�cA�%��eO���ǒg ��Ӂg�����U��մ�*�^U,�3g�{i��b�[����CvR3)��,��r{��i�S��'2�'�Q���R�>��j߻]��
���9((�=7�g�'�¾�V���BJ`^���#�J	-$Xy���	8S�wM��d�0��z�K��}�d+S��}xd�&��mH���@�0.�6�-ǭ��5�1G-,g@��s�boF��g��.����*D��+�A��P:�a�״f.��f���i0�!����J4�BM����JZ��)��?Ի� >f1ev���؜	R��؅l'=JD�6�lFnT��`�oщv#Y"#em�>���ə�*�
��UM_�_�2�pSC�Sx0��*68�]54_��� ��T�V����V���:�>���&L_�Ru��0�,�Ϩb����k�Բ�u�w-���X���Q���l�?T��S�bQ1#.�u�m���@�T����|�9��7v�ޣ2�P	���_X�/�R�j"�O��Q�����A�k�	)i�gR���]
�%?L�{��g���v�x����ZT�!5�%+��ɿ8�Z�~��"E�UW��$ ��+ʊ1�tw�X '�A�=�b�B�Uٌ���xl.a������|0	���	��G/S"kCax@��8�*�c���C|��	�z��7�7����� .�M����׽/w.�}�$���U�y)��>��US�PV�js��qe�dy��yo��<���L��F��E��|Yj<Z�b�z���0o*��O�Ƀ�4P;�v)�֒r��FTIw��y#�s2�6�N���"c��]ψy#ɟ���b���٢/"�l���۸����IS�0����a:?��B&)bl�M�<��pT?G=)Z���#����Ŷ��4ۍ�l;tXW~L�/7��볝�ϩ��t��_�"c; �������«�_~�_#�k��&+���>Be+�o�!mX�rX���x��hޔu)���2�B��H�ĭ�g�uë����j`��R�X+m��צ[�ւVǫ��:<�p���gtU_�(䋎��pP����}nMIj��?��L�A��n�?85�2�?�#��WQ1:��C&1�28j$�{tx�%&��\�8fvW�<�)$�S����:������?��S�h��#mx%�s���W��9�K�w�j���m�*�� J2R��vx!��!]���#敗�緵�Ƿ�����}W��o�!�#�x��/$�eX�-{H"�UܯAJh���<��hEq��;��OA~�]��0��ĢB'$9��j1��h}d��8���3���šg�:�c��W��[�A�$����}��]�����d��_?��"�o��O�y[�C�0�������Q���+�^ppMu`��7� hH��������������+����J�ץ!����M��'��H��S��?Kϐǻ���gI�1�kՋ���B�b�u�8�4R݈q����#HM75��Z���M7w��F�5���͌Q��^r��׫	�m�v�i���93�Ot���_��.��ٟ��.����8W��[�ǘ��(W�Df
��R�Ո�gL"C��v+�Iv���Ý�x"�{H;��l��9����R���`��ߩ�N��y|o^��ؓ�EҪ:�+�#��ɶ�
��*�K��Q;��8�1x��YU��B^¹���yR�a�BA��/o9��MqxW���>�@}:T	E��M��n�&��V:���g�_l�|0Q��m*�n�&���2���mSeR�&�cx�z����	���6�Tx�S��i��=���?������O
�bc��0�\8���L�"�ˋ�n3���t�O�,H�e�H@~W}͏��P��V�+�T`xr)�TOLb����T\���1 HWQ��ʃ}��ԫ�ŝx�1����y?|'x��.���٨�+�P���z1.�����>*L�,쯅�$~��"]O��N$���p��u����"NF5{�Q�m�O������MI����j�d>�u$9��|g� �h	�}����,-�\m���\ѦqV���M����/���7n'J)��Ts�w!�S�5��aE���\Yr��*�<�'O11�Pc&��ߜ�
K����Ǝ~��NB������Q�����@uf[߿�W.�`���Z�⤀�L$:����m��O���|o��{Ԣ�""8ȃi�M���á���wm������c����䚩��;�tr�e�Į��T�q���6I'� �4�u����2 W�rY rSin�����_9E0���4J���	v�'\5��N�ˠ�*�3(�� �Tߵq7F����B�'^-��3��������ej��RSv� ��>���o�M#1���|#.xmon��0=�3F��:�PE&��^BM~�������T7�&�fWr/9/�1�m������e�`YK� �.�k���0��]�+�#0a��V2�ZBh����#�cO��U���#!N�`¨�Tu������]Sܽ��K]Y��#�7�?N$��?����W�IT&Ҡ��63�j�yn)���$}�><熶u�ߚ���T��.���;7!U�
c90\��mx�.IM-�g��k1��w�v��7e�[��TL:�����!�+:��i3���8`�f��M&�VH 3�[�d��$}̯�"�, ��#w�ϔ�?�bcqo�)�QL�6�2��3���jԂ?�vk�i֦��ja�IM��qb������(�$P�N���Ŧ�J�w��M5�-p����?�Wd�C�o*����ȝ%��3�TjJ��f|5�m��,�T�w+X|x� W7���*�C����N.�8
T4��}�T��	����6�+yg����f�z��T�/���*F-zj��&sU��/��3I,/��)v!�|�ĺ�t�=�47�bj����k��4wv�H[9<�1�ރm/<�R`���T`S��c����b�3�����L��4�	5-��D��� �e�w+z=��	�N%!���N����j��%�r��O>N���8?�)��I,?3�d����K��j��J#�<4�b�h���L~��S
��\��v��
-/<=`4��i��7<l�*ڨ"R�,�r�UFU���n#Ü���k��;�D<��A�����j��} e\@��Ж�R�����Sh�lzU ��t�jv�ۓS&'�V���d.�	0��ߋ�o���}�H�c��ešA���i�U�����C?O'�ԑ�Lp������r+�P��5b3��g��zz���5~b���`���q���I9q�}
l��J0�L�r]E�1�c��᪓��?�=��o�OzU��s£�NG�v1\D"6E:���a�^X����D5hU��W��L��s�DV`�0�r��-p�g1�H{�@��]t���T�� 2U����5(gd@����K�*iL\}G�"����pQ�2l��+}&�Z���9lݠ���ʑD�|�Uҁ��[bed��Q��Y{ű<O �FU�:��	�?���c?��T��*�h�,I�@$7�'�eɪ�$�XL5H�����2	h�8��?n����o���Lf(�o��0�i�8�pK�^�����ȑ��sa$�B�;�?s�*A⃗�,����ݓV@څ[�(�!��wJ��|ğ����3���o�6Y�e��&���cp}��~�#����?ҵ�"�&�*��fETО}��tխ�Dq�Se!=��M2[ĉ�����k��]��y��64�Y뱱�p����������3��A��f&�\�$J�YOW_]��#��ʏ�t�)�s��3}�-��eHM�]�?�-��fkOn�M�J09���J�i9*���Y%�"��䵂ڙ�w��@wf�A|��x����j�H�rn�j[*�q�l���#jzS�B_��U���T,w��`�OM�ٻN��pC�C���	I:�*�,b���:Y� �C��<��PQV�=a��|'�<�B��.e�����a%�i��2w��]o���>�{�S��u�3�1�Nc���){��把g7�p���̑�	�B������Kc�����2�ʵ��v��[��'vz�#Ó���}8DÚ�k�z�1�ᰐ����Yko#nc��L���I���%�����h�v�B,5X���%���T:Ɗ���H�u�����p������!��r%H��c}�x`s�h|���ߓ��\*ɰ���Jl+��c�@
�|�z��f���-�&��]�i[L�!���`	���q�yrb��㘰�Q�C::����r���l*�!%geЧ5�f��O�=�;�mC�ެ����S_M�J2�����(�k�#�Ō���t�3�%��e�WG��
<�W��_U�s������c�k�.�)��'m���n`0��U���i`���/Nmp{?��g��no�t��\� Ǩ�F0����x�B8�O�B7;!&Nx3���1��
��>�U7�R�K�����R5��w��~>�%_��`�G���(z�m/-��pC@%��ij�H����$�E��OFH4Xj�J���A$���k~$�e�}&|3.�G��ʺ5?d_�{��z� �<����z$�\-�si)s�`v6_C�p���]^-8��h��yzv��{�[e��aq}���:�wvgW��m~�?l�do���ZN�]�ϝ/}�x�����ڵdM�m%�H:�7ܵq)h�MVk�>�{��t꽼�\"s.(%WLjU�j�֥VW�e@�K�9ޙ}��'�	f�|���-����͍���(�Z�s(�r�ӼA�D�����56v��9Ͻ�YMڈ�-@h��=�(K��$|!����]ܗ�ά����n&Ґ�`�I��~R��I3�ý�j�'^N��,��E���ƞ�I(����	"��� ??�����v8	-81�/�̎M�sj�,p�.���d���O��亜�D8f�����fM� O,�� �GAUϓ���4�2�0:���b�`�q��]O���]�Y��`� �E8�{��S��Yy5��l��e�)Q�I�։���3��+�b�{�����3��fx`lltY/�A���������zW�w~�Y=hn:��፛?�b~d<��:��S��u3U�m�U��G���������A��h�� +�~��*�F��4 ����J5'!������ta������yn�
e
�0��62�W?t�oQ.ѱV@Vn,?*+�c	�s��T)i	�����"P �{�-ݜ�c5e��F��{Z��mﻡ���
���ۀ L;L:O���}b���oa���{j�ߝ� ����dtB���eѼn7��pM�5�����{���Hd���l(��`�A��LBQMD�F|�iw���i��-�b]��͂��p��P�nY@���cT_�.Ywo�������jID�bh�y�Q((��}����h���}��� !Gۈ@�ȁV���C�p�0πɽմ��j��{�[�Ht�m4oJ lŘ�Ǽ�T�?�*^[de%y>ɐdS;&�'M�����t �W/ט~R�~�k��%�؛̓BDT�l{U�<�[��%�����i_ߩl
��B��E����zi8=kY�v��$�K���|ۙ#2���dɳ��i����@���;��� [L3À
��&��ۆt��5%�e����c�~ N<T�9y�Vo=+X��Ei���g#���\�d�9��Čp3�ݦp}e�3��>}Zy�N��z2f�m�c�~��aF�>KȌ��;�Κ�̘ؼ����c`H�ҙ8d��	������e����x�#�l�C`6�Ҟ���mWge���Z�CPu>ts���R�%��Ȧc��]�W��==��k��0X[=׮ߓ��N�|��+�^b ���o�Z_G)�3W��j�92�l{(詭��y:����n<���&{M��acpxHBE� �P*�&�����gO����q�%9D�Σ��
^:�1���,e?���LwCM][��iwD�v1<r53�$u>��BU�ҿ��_'�$\�R5�9�v5�7;}w;�m {���[���G{��nD��-���l�^6�:nj��ã��7�=��[�݈��ib�IERCٱJO�&�۩�.�4�-H&?��7RK�-����w�Ԓ�c�����(B��̯"��
�������Aۙ�0��먝���gdЊo�	�˪��U����z�·����c� �_\�k���c�-�2VpC��e
zo0�����1Ds����s^��Og:��f�h/�[��xU6���#���޼��ɞD�-'/H�\��a�l���}I� �G&�j�t�sK��g�bW��\#�=�� ei�΍��4���� Ʋ����VI(����u�f.	����I�����k}���ʅ��-�v�:��I�Ѯ����<����x�=�鰘#�����l���6�js���T�i�N"��W{��j�h��+�ox��̻ C���)ѓs�E�pzx�͝]��q��J��͙��{j�a���j��+��l"��΄.��+�[��9��s�*����P���]��z�s���fu�t��'�ZY�5��/4m>��$�.ӎ��`���{'�ǋY~V�R؛�(��O&}��g����N���ڐ/6�v=f��(9Tl�rXQ��� }B>�9�6b�sd@%��� B���y2W=�.^�^Þb&�^ԫ���Y��ؗ"�h�ܪf7�I����d��l֕��t���?�3��8S�����Y�󭆊��x�^pNJ����1��Yǂ���1�:s~�������@�����h�a�b��%�zh�a2��hOzfl���G�e��ӟ�e&�58��Z� R%v����-���$�O�_T��s�M�e�>�{���{��Q�7��h�9 �>..*✕=�[j&d�7bz\x��P��r$�Y������Ck�7ڌ��>uK��d��|�6�ǯ���������q��L����9Z����q�j[��6�.BZ6�_��\�� 0�콳6�������;�|�J������}y̞ޜ���ޟ����t
����Vj��'a�׈�BW����=�@|k9�4�W�G�,q��n��~ӺM@���~}v�EY�΁@�U����B��ŭ�AY��―��=�Ps}��V�m�E�3�����H@�����S~~˄�4��|u�խ��-�����Q7�L�fTE\�|9������� �*˻N�@�)��
�|�+˔��x���P�M���\��������6Na;���ĵ@$b���d��q�7n}��1�^���cBW�y�=�_�^絶����*���q������� ��ǣ�]x�� �҉��Z�>kN����2V��%z��d�t�󅹌���Y�ـd��<؍//�Z���A���v;�>-fUy���yz+��ܾo��sK3*���/�&Z<6�S4:�s�U�V;�����<�J(&MF�'_��n�&׋�ʭ@��?i6�������nk 2�֤�b3�>��
\P�\�=~������>�DG;X���O{E>_ �
�UV��@j�m�A�����p7-�������GY�q��^
���?�n/�\Q��Y���ڒ���|i�"C����/� k�C�6" 
���9�N򕡕	�8��IZ�x�iO��G��0gD���
@ț��޷@����^h����B�o���v����S&����!h�]�" �4i ,[ϐ�����{Y�qc�&[BA�2X��8�x{�!<H�'�zά�G
 4�;�r����� 5ҷϘ�4��j<y$�ueB�w��P�ԍ�p!&���ߓ�<Jb��^��R�ޏ'l��P��h�-'-�)�8]M �L4���ͬ
��?u�b+��q���o�̑-nAy�K#5S�a,�ˁD���鱃7Y��[�=��Lޯ��ָ��h���L����ۑ&q�}�[݄ɞ�Qvv<T��n^��&JF|�r����H�����Wr�;�h|��"}EH"r&�0H4�L~\����
��.�E,��v�_<��9�B�Q�8����J_~%�P�n�h��l��e�����gN�,ը�
�����.��w�����5&s~��P�P1{�7^�D�v�����P)����C$�������:R�6z5$<��!�~$�����h���[S��y���Upm�JI\��k�6�f��A�Ɵ���vF<�?��;�q7L�]�M�1��b�R������ŝk��V3���WR/旘��Ɍ`�jQ��J:�t�$A��[�8�=��<����Dc�z4:���O�P���t�/�>�.�ߜJ�ޕ�:��1�d
�i�a�,�����3�7�8jH{�,��.��=�v�GY�-{�ޏ���~n��5��ΠMN �4��z1=o���m�ZG�.�l�An�[������`�!v��� t�0P޶y������{|;n�
v�E~#�����-���4��[�?IO\�X��t��S�����\p��oHa�t5�b-Էd�u��U�:"�4�>�t0'�Glǭp����<���r-�چ�p4}�<a!��a�|yFu|��K��N��z�  ��n����>:Z�ĥ���b�M9����BL�\�������#�~ �i]���]8�ݏ�:r{��y�eN`f3{#ާ+���k!����U&�Lа}Z·:�5?Q0HqÞ#ޗ�o!�]FU��8�5��w�TqKq_}�	c	I�|R�D��&��_�l৕/���Om��w;d��0�wfKb�����y�(�(u��\��u���Fa�������L�A�\�_��jP�bPihX����k�!��I�y�eA�9�f[j�3%�_����M�T?u�>��ru���c}/:Bz��Q��υ3��=�4�d�g��0&��?�>m���FȌ2[b���6��6`���(����^8��#���l������۬��&__d�s��_��ӎ�٘*���oI��8M��,����i$�5#�#�� �c��,��|A����2Oӟ�&�'�6��,s���z�����/;�G���.�Y-d�}VHYݍ�Pg�Id+q�Q
�}���3��J2��F:弜�z;�yVU��������.g>�u���@�;r���L����,�ɣ�DԏM�Z;��F��J�IXb���cS��ɍ7�*�RX������+�X��Y�_��a����������|xg��q�7�u�c�~C�eY����C
�]@҄7��p�5�4���]}��lɑ��
yv�\GG?��fz~��*�Ts��x�
���u�]�k�W��Fч�	�Q�������W��׷h+��M�hftK�3<���S����7��|!��~�y����bIc� �v�w��cb�����S�J������Q�������X�Сň��XI��퇇$�߼H���~� P(u��q�������T�L����9�dm�ë|fUr:Q�QX+d�^d$���B����QX)�q�G�+rrr�J��x��u/�}[��!iD���[���KQmt"�Xͣ|��5��]���~�^nc�u��l��c0J�o<�C�����E�k~	�o0嚱{E�>�L�Dp*:j0��_LE>�Fq�o�S��fKگV��ގ��yk����銀޷d,' ���!�
m�37�^�4�1��8;��]rfd�:̌X2�bo	u�H����E�C ����&�2�2�W�uE�J]��\i)I�av�|=#�Z���ݬF���1��Vxh8��{�l������ޘ���������p�����f��_�l�� ���znl���A��C�2&�V���7+��!����f���9\��M{����-����>D�"��[=Ku�@5�i�H���7�8L����:�۶0���/.��3:���fޓ�T�D��b�e��[���~\��S����%@�����͔!"����G%����$z�)bw&�v��'ۆ��7�i	�M�T���"����c��jD������LF�F��
�!�4�[t���͐�wFd�o�T6��s���~���f�Q�I�s�����M�
L	i�G�Gٿ�T��'��ʴ��~r��ƟLw\�)����\uN�@���G���M�s���	�̥�M������[M	]\Y��U��d�2�a��$qv�� �<ǁݑ��
hV�o��(H#^X�@T�d��kl��ZW\G���\�D���Q�>6
Ѣe|ǈ�R|Ȃiߓ�_�Y]>�h/��I.��ՙ>�p�g%�-�5 ����g_���&Uӿ�4�(�zs�A؄���ɉ�Vpj�E1���x3�p%1����鈯��vBʅ��F&U(\w��|6a��IhDI|��[�1Z��D��i��q��}]��ߝ,�T�y���ݾy�*�7�*��n�F@�������<���ε�*�22��$~��T��h�s�&]E�Vo(������{}��
��o_H��.O�] k����DhF?�n�YRq8�(vn����0?����`��ƅ�"o�̥��cx���E�Z]���l����@.dd�)M�c���D�L�k/�\�>"Qa��K?6|��q����ff�i�y��XC���Ijq���>�Sg~��hr����ř�N�f٫	ܛ�ݲ��~�1�#��p$�yؾȵ�s�����d5q�=�,���t���iyN��Nj��tL�/�ﶵ���ɉ�e'�����vn�,�·�_Y��s|���~���t���{n0�c�����ŢR:����݂w<L��*�i��\��t~'�>Y��f�aPꔴ^*Uk!��|4�����@�v��A?G
h �����ͣ51���/x�3�I��h�_����7�*V+t��]����F�v�:OLM�}e�$�����Fv.�͒�O�R�<���u�F��㖩��?���h�6.��"���vkR��5�JYhh�5E�W�6Z^���[��)�	�_~���3CB=��9�(5���������� ]<g���������v��8U˕�Ӵ��{�nӺ��o}���
�o5��a���� 2�]�E���5P��cl�n���S�6_!V�}�#��bi�j�h��Vԋ�Qo��8�0㓲��._n���7��aD����C��1���ɱfM7n��k��;].j�k���#2 4q��7ȃ�̝2gM���%�G}3o�C&³j���b����I�Jb�MkZ�i ~ g�>e(�����������ҙ�7/C�Yd�~Z(5�7Ii醆D�*�A����]��X%9�E�Q���w�[�q�WST�A%+�-��/t�b��I��������^�8��X���L�{���EX����`�>�1Y��$���? 8�M��gP�����{�#���"/h���NYn����7�W�$hu�z�KN�B��N��� Ѐ��,l���f�b����gkV��5ӟ4���O�pG��ø��s#�����>����.w|��Q�LBR7:���O�Mݽ)]o������k���s"�ΰ|1:��f2O^�����H4u�zGN_���p�����Z�^�?�x�b��������v��`�<�h]$�89��o����sf�
��2|�S�zE�����e$/p���`��g	�s�0R�ĳ�{q��Ӡ���,NA�����ޯ֓e.uǹ��*����{���_K���qG	�2���eT#��|��Q��N� �3��C�Ņ����[S���hi*��8��L�
e��R���T����sV��3����j�$m�`g�Veۺ��v�R?�<����C[�5x%���`ۊ�pq���"ph����in�/'�t����{0>�����AZ�V���L� d+�4eO��lԨ#��^"��܏�ZK�7�G4�����.5x�Ά5��b}ꁋE��`ShQgͨ���-j�&��v�`VC�+���J��z��9���"�� h��F��Ӷ��D)亢�3�q�$<݀�5D�x!"w
>��+�.�H;�h��/�����{oCۺ-U�縯�q]XX��Rk ����k�ފ�������D �`���.�x����m�%��x	��>�["���y�ǲ��LW*�I4���I��!��)f�� ��G�m@ze	��(ح)��tX��n�cNy��Ǎ4]�?��sH��E �#V��t�Jr��z�/b	b��c�B��;��w���$s=�~s��*U��Sc�����!i�5�����2�;���^.ߏP�Nz�yE��ゞ��=[�9$��y+�y>}7,�mw@^ͼg�����~{����������>xT�ݺ��#15��1�߃K$cv�"�q��O���zn�~�������v�/b}�3H{��]�N%�{5�}������4'ec�L�H+�8�����!u*���)��_�NM6[`!-c�FW_ 
>wH�n>��Xƴ�j��3A&<��CI�G����7 
��D�+:��~�p� �=���,���={��[����0�%N�|���Jj�O< �I�\'V<r��(�p�z���&~��S�e��N���*�xo�*�ǉ�wg5� {�ۏ�'�|�d�.�sc�q�Ƿl�����j���EAT�D���R�w��+H�5� *ED@A@z�%�BT��tBh��Jh���A�s�c�W�=��R�^k�������=�,��jG�Sen��S �ۻ,�K��3�N��|N�!|,�|$�ΜcB�褎wI�7�i�$E/(	��q���������U/����l��mM�˕i���r�)�H!����]ߡ,�-R�P�{�{��{��k�ec�d�4:���Z�~��?����G� �0�Re���d�
߬�SE�#��G��L�X�W��3y��Nڒ^�P&؞y��/D�L]W��ȣn�>H֦���aF񎩯/qB�	h�:�?K���U�O�g���.�nkH�����³�;*�2�3��a�!��G�`8e�5�)�-��q�������u#
��I��`�y�:����t�)Q!��S��N���k�5Ғ=Y]%>r�F����=�q�\��l��h Z����% ��@�I�]���!����	��"���!�6�@ڵ��@w���7�_�C:�M�&��-KFPf�1��!�n� =�A�ۋ�ҋ��Wyy��ӛ�p����5��I��8 ����!�D�����[Op������\���S��P��@���k_zE��I�n~�1]��lI*L~� ���R������BZ�x���p��>v�&�����ʒ���R��K��-�~�D�b�� '�<9��?��E��:'�o�����}��H�N�C�>}{J�F�iL��9��  p�Z�G���^m�J6�ӏ�e����؊�zb�4_�2������G*�.s�����}��0إ@�$��;����*ʎ<&d�g����[Q �lK��'^b�Wb�h�n0]�<�����e4���O{�:�^���I�J��5X�M@�GV��}��G��c����Z�����ѝ�N��BZ����B�	�|�R(q+z+��F+}ނ�M�jaQ�d��U�|^��g?���6��z��Y���מ�M��<�� 1h[��xu����e`����)BH�$��٘F�r1n���)/�=�qu%XC�+^2߭�R��v3K�1Cu>�=��J;Mͻ��Q����ܹ=��)Q�\�!v���SE�ξ#�gs����R�T�k��}-�i�3_�n7��)T��B�2���=N�뒼���Pza]v�m��ۛx%������/�o_�Rpd��X�ʞs{��@B��ok���N�:�J�}����Cx&�|��5J�qN�) 4�P�W�����[@��(�>WD(jd��.�)t$���Y��T��3�)%|��b������
�>MFq�=U�>~wŤ���1�\AZ(B���_�O
��x����ܰ�i�WPT��n�s�ܴ��#n�Q����!�n��۩xܔ�%�gT��Ǘ��s���H-ҫ�Tgʲ>.O����Q�a���VC=x�{�T�5�jc\��ٍ��X�-
��-[N�6x�ΕbeHvs����A��8-���	e�k����f	����\cD���P�*�:�=.fT�޺k!m�
�F��-l}�W��~��	���Y��#[�ߏ<b���ŉ/	�Emmԛ��&���ў��eԨ|��)�r�_�A��b�a�-RSkH(�	�GB�cas1�A;���U~�0���utr?�\^lK'�`C��wi�\�&���{�dAc��*S?�9����f�w��,J����^>:��,l!�8yC��<w=������))3zњ��:�l�s��:0��ycm��cB�5|����<���7k���b�ל؂�.RK}�?}�]V�����kr�����9��}���d�TT0\��x5�k�g��c2I�ӽۋKK��gU?������\Ն������*�Ŏ^��r$�zq
7vt�UyoF#�RR�wM����I����{��A�C���h��a�J�[��":e�����=8���T���?8��2%���������'r�ˋf�BZ3��BZY�h}�|
��&8�>S�.�o�ͻ���O��'������m}5�c�;X3���m�zb��9J��2R��o�����|% d�xq���_^��y������{��^�'ĿxBxI�⛇2���H�L/>���#y�����jh�~���%�z�i��$�j+�'�פi��c����N�io2j��yCM�y�)&A��|�U���U�~RH�cF�����=$U��A�����$	�����!�ǏWu5�_D�{��F��Ab�8�t����1�1�]�������s�2N����J&�B����'��4-e�*~~�וh4dF�k8SV�֖.oe��~$���v$T��O�/�R��뵠��gМ�:t�JE�Kŏ�c=�&E��i�LaZJJ�������~~Mj�"Y�)Bʱk#%�D$�?+���PX	"I���O��L���&��&�˙6V���1�k���_RR������������G?����=9�cb���ϰ�������y`���ڴL�~�q���}��Xf\mԸ�Sk�����  ���`z積1�=i��^��,,}�Si\�OĬ%RhR�t0�������w$���6J��PEͧ����'����V������X�ii���҇z�'��nP\����*�����3�����Cf�����9�S����k�����;݂�P-���4��O�'8R���Ƿtgc��ua~s�zo�^�ώ���djr%���au�gm�O�jZx`�^�˼����^��n�TD%Eȱp����g��(ی	+/���܄�h�m}��<�J�K����0�d�{L^vo��|؃�6d6�F��ϣ�����N=��ᾒ�;�F�$'����*�ǹ�a�G�5*
� �&�^i�Y���;9�>����4� �t������U	�G���/J��P���b�?��΍'�^�lPT���xM'{�?�ka����%�{.S�'[E��Z��ۛ�cy+L��ʵ�2��y�Q��ڇI�ݶzm���B��Q�Mo�X��՞�Rl����%竤b��;����0�%���	���;�̝�Ȗ~�e&���/���L|�^h'��ш�q�y�3|�1�  iX�z��\; L1 �e�̩ķ���71��qx��C&��_�,��wML����'���k?��ܨ�zb��J�C�p�C�|��#��>�8o�l�d��P�YF��wMsҞ=��h4!є�bY��棯�^X2�'m���a��dK�n�NJկO��t��ĝ�QKL��t���+��#�����"�7��\�L��%�� ��J=d��	�޽�@����Dp��14��B�>����_"�DMnWҋ�*���@���k��N&#�ʈ[�ѿxp>]��f2�)���DY}e�3��2)zQ��x"Ϟ����&@>խ^*�]L�TPX�ſ���~�w��łR�Wo���'�v�%�=�)b�׬ H���8����Q��j�"�;
�a]���nP\bb�EL��:WȲ\6Xy�f�T�"c���{�/
���������g�=b-YZ��ؓUX.��>��T��U:!��x�f9���DHL��6��)����Ʈ�:"����F.%jp�IG�d��R�&����a\z%�~e�u-�!����)�7�Xa�JGW$����e�P��&�FGǎ^��,+�R*$��Fo� �~�	f��J���<~�M�vd{E�իW�7���Ĝ�솬w���D\�1$T�	�L?~��)J�F{�1~��O�Z+T��j&�@yR��ro�G��臥�J�d
�j�ڗ��L�NTք���0 |�Z��H>���=P�"-����\*�U�k����;����N*6�P]d��ؙ�c�Qd�`�9;� �[�Q�֐u��S��O;%N�5�B�+[��Qʤ�� ��}\�yU�����s����Z�ms���cx���"g��3
O��t8'����@x���
y5��v��g2��Z��s�A�+z=��`�6�Jۮ(������I~��%H����>�/u(��Ih��ܴ)���>E���r��7�f�7�M4��3D4%�����5���)錬�L��?*���u-��q�"/�oF�v�<ο���\���Ԩ{8�E�����)&��*K;�����@�l�)���_�6��܌p?���.�H��0�}o_�'�������Pɋ�����j}$,ژ��_����n���G.Zݽ�&�s^X�ouР��855U9jy~=�F�yV�b��z��տ���zl�a����1k�[��k�ɩq\��U��߼�R�9?��df%�����5��uf�իWB�➞�x���#<k8���8e%%=�0����p4Z�:�B{�5?l���$'�[�&j��;��!i?��^���H$M��p	����A*T�â҈Q�mT�z|��GpW��L%����N�y'��͚'Tu���oJo��)�=:�C���Lׇ���M���,>4����~!����٨r@�@����|��}��?3=r�����/�����dYe�|�ʓ��C�O��	��������Ǡ����6�vj��㗷�5�{��Ւ؋�I-#L2A�ɡyMPr�gFщ��Pr���ʶ�ӂ�d��������?�N�!W��""��x�O �^&���|�v�J<�u�l�r��F9C��#����g|�M�۵�#�:��M����/���|d�����LÌ�|o�krW�w���z��>�:\����Nx;�TV�8�@<~�,�y|o?v�GF��������U����'�ċ]�Q���>3� 3���7�@�o��̟���D��Eb��ŕ7g��>D���@@P��X����E��`�V����ʛ6������63����C�7�cf@C�jt2՝#p��X ��x7ٳ~c7��1��W?��r16ˆ���3o�?�m�ZKL��*�����U��{ITm1b+����k���]|���Sp�� ��~�9�ؾ\�׌g0�������;�%����	g�UE��f�X��7��}�k`8��z%��ǧ�����r�rm���ݹ�oy��/�V+8�G�F}-7�0��~�;� ߯�V|a��4�+�z����X��M�'�c d|��[8�M�/��2�� Zெ���RN���Cq�!�/�<=Q4���.d�qOqv��+�>�_���>��R>�D~�$���1�GE,h��MP�����O��wl1���Z�3�i�� � f������V����y�?z�Z�U��\h��т�r�f7e�������u���q�[�5���O	W^^��a-�X�V�A*?�^q$.&F�3n�Vl-����d���#Q6�N��1�he�g�7�ǅQO�q���NЀ8��Y�;���69�n��z�ZQ>���!́G:^/���5�J�~nz��H|f3�mw޴��dSP|zc���KZ��m/����V����C��Z��A�b@@3	e���7"NɎ�J�˅��5�:�f_��߹Ɲ��5�w|��Jf�bW'Y�9ب�'�εz'����PΏ�z�d��74YM�*�:�܋�GG��"��+��mx2{��P�\̤�&H�4�"KS=�Ye�;�CIE6��ƴ���ҵ(D��C��H��JM+�e��:��+xݦX��9OL����"-f��@gBO?P�$����o0��"���������u���-)��wPi�ym�OТ���E%�Oa�p`A8>��	A�	~��7��P(�N�W�A�z�71�=��`6X�w2�f�BO��*	���Ϩֻ���]y#%.� ���VH�g��>,�|,V�uU� �[���P�_�eL�_��Cv^�h>�&z+��C#o)&�\[:o�3�6յ[XR����7:�5�=�ES��'�?[��`�Y���ܻ/����������g6 �52zL���^[��i�SW _�ݞ�O<���32?�8�p�&��D�&�щ�|j�scrv{@������QL���y�@Cu��G����ϿJ�/���o�)o�Y����>r����d���9�1�>�v��� j�����'�1�I��B3��Z;�?��@���m\�>����~J���%S1$���H3O���Z���#r�j��5*
��� w����V�.@�m����HVO����s�'�x��y{���=^r��Gj�U�G�"��}��Vv_I
�B��T�iv�����V�kQ��l�?E��i�[��QM0"�����1��̬�{3ѧ�\OaI�dl�$J�0��k���'B�a�' 4��))�)���]�X�)��w�߲��ON�|�@��?��Ly8C$IM�T�c1x|�3 �K5Q/[��N�����{��<v�%�uq�]]�o�܀���++�q�~$\~#!)����cO���홠�m)ҧҝWؿf�"B��6k��P��րχ�1��Wi͟�o]����-� ^ׂ=HT�2���^Ȗ�U������˼��ݰ�-.|l�=/�(59z�oJ���pY�ބ��������o]�(ص'3��ֺ����}�IB�RJ�Ѣ���52`zhH�TL�H��~�A�d��4�+t��+ی	XմT���B���[��\���cn�+u��mqwW��R���.��M�zg��4� �E��'�����l��Mtm~P�G�+����v���L��=�a}[����	SN���c�/��#�ӊ�y9����[-^�'�B�c�rNVc����xM[��%��!���.�7��3S���ӥtr	�����&#��=>VK\%���T����ƞ�w���W핖�E���P`�zHUȗ��!qK�C�(f7�Х߮+���9�a{?�B.��Т�@ѐ����U�2����uv*n�T���gJ��)��,�Σ�3,׸�2��;�ds�V�_>����`J�������w�7�j�e���>,�z�����+���N��4�(�z��I]f�S ������r�ʽ	쉶�i��]�i�댲�����rϙo�=�m�e�&#h���|�|�$�B}u&K�� ��٧B�뽖��'9u���ڕ#��s��r���]ɓ�����>"j�NQQS���Ŗ'K�V澷���tI�kv|�(>C������%$'��Sꞡ����J󐇛�z�N�	Ʊ�<K�ڼs����3N�'v������ַ����^�Y i�����H�`�����G�b�k:�:��}����\�"@�]�z�iM1�mH4��3�!��,k�Ԉ����b�_ִ��+�<7?�XCtޤ�ω0�5.��l"x�F��C�C���Lm�X̢���2w�8���i��^��>֬a6z-b�R8��d�gZ��Z��z���Q�jH��5���v8镳2ښj��֋RR�M����ץ��J�yp¶�{֮�^�b �.���7 ���O=�t����D��F��5b0G�$���y|�ܠ.-��U}����Y�[¨G��Y�bHz��K��f?M5�Y\��K��f'�������j�q p��C��H��v��K��j�6�Q��C�f��qP��Sm�d,�.�:ʘXs�F ���;�ؒ��ҽt��L�����)�M���6[��h�ëۿ���,\��c_��l.<�?�N�<��̃Tb�1�ǒ����ɂ�q1/���J䱇��tͻ�{�>c��Xr�X$˝ӌo7/on	�7[�� ߫����x��8�@��ZѷOƸ'�l7��`vR��G�P�5@f@��2�D�'6��X0�m�"O���R=Ǿe��R>:i�5�|\�r�%C���LY���y����m�-S[�V^e�*s-���_�j�f�Dآ8{B�˶���T��ĪϷZZO��k����]��M��*��� �wl��nc����5�JO������$����6�(�M+z�҂V�";���Ϡ��W�p/�d�?/�R
��ʿ��^�pH��+��*���5zd6K�	��iRe8�$l�Y�pD�O��"p#�|��CA����#T��1�C�)V��(1��Z7�upߙe��Ρ
Ł��1�o�shP����p�Gkmkjzm�z�����6��V�������5��:�3��j0���G!�1�����Ă����>�����V��������BN���K�C9�F�CS��j'�YD�����=U��z�*�o��f���.�[B�9L�~�#7�#���:�ܽu��Sr)���go���w���h�v�V�)xsʿfr�P���u�#O��v��5(��G�4~[ЪK�҄�T��xu�E�wWM��|6�R fs��)"�E�c�֏���_�Y[/�4&�|)ryef�޴��L�=d�`��A��=X�b�M6�W'>�n�>j64���P��@}�L��&��!�%t���
�}�����_C�Nq��q]G�T�G���{f��l	�b"��jc�Z籟�R'6��&|���>)*�zJ=��p/Ȩ�7���fKve���L�"�r������<.�Z{��ؑ�IR���A���>l��������6�% �r'����6�F�Lw�gm��<8=SQT�ez��\���QY���u/�Y�>;^��\Y��<�Vd^������4��*@�<u�4�[��	��U�1Z�pĺ��b�N)2uXF�]3e��Hm��=(��V/�f�n-ߔ��������n��6��:�r:����]ss�ޯ�o\m�'"OM{{�U��#����~!���t��%#�>�&�涘 �"��%�ٞ�������IZW�o@�_���XԹ�x� �1	�׹�ܼ��!���N; �*��A�>�j�B�<�9zۦ����+ut�>ɘ
۽o�-��q�����*�Dŷ�b��@+��)��K��y�[�/GQ׈WRS���x#�Ej��Z��㏻�����r��]Ex"#�"*�S�N�-�Ddk��g�#j�Ï��P���s���\�-���˴'ּ��tЇk/0���6�U��eA��>�s���?�9*�ϡ���;rh�.jz�{n���,�#�|��l�c5	A�o�
������67���e������7�p�	Uz�2;��I���,Y�=\WO�YEc�ײ�ȥ�C'4��X(��f��k�dT�E)��:r�i�nX�V��^�s�Q�����Hl=q�wz=Qk�t�
�z�P>�EA���:+�U��a�о�}��ﰠ���-�@$�����\��<9��%�$�s
��+���P��,�R�ʝ2\��0�}�J�f��Ipꨣ7��x�@�؉Y�������g�o߰��ի�S��hV��Y��=bZ�{�i�t�&F�K�/�u���t�3&��\b����V���W�fN8z�$C������#~͓�\��

O�~���<E/]	DY��P�<���d8i�H�|E���m��-A6唦Ӻz�^w��y0.��@�~��5h�`�@���VՍ��/�/6R博�����y׋x��#�3 ��͌���Vz�����#�}���4;�!c�R�TD)�.����	��-aL�g�^= "�y[��I	�Ҝy(+�z����d�Cl{Ֆ�F(�/_�7;r4M���$$��3h���1��L<u˧(t�oe@��a���ٝ��MZ�F��A�
ݗ�{�R�W�X}Ƙg�j��R�u��k�1M�A�ޯ�0_?Øz!1c�V�"���v)��?z0������oЀ?l00���'R�mҔ5H[���*`�~��>lv4G�1q�7L�叙(v����3_�o���u|��?~t,ț}C_, �sG핻��g\,ʎ��s�ؗ�8��p�r��&o��2/�u��'���o�q�T:zY��f�_��c���kN�V(��ijT�5��'�"4 Q��*���\�l�B�y6�^��#EV�H¯j�����g�Y՞���U��;����\��<�����]'q����yĩ����݌gsq�(�`�J���qM�MI,�h�N�ؗnD�Y�ln^��(�i�����PBXX݃\���b9����I��ӫ|$׶K&�3�\ba����#e*��7Vk*-5m2 +��}����fc>����U*f`6Y�"����)��6�Z
툅ו��/T0�0��>G:	z7h08%�Զ�)?�r���{�S	j��LM� 4?HW���`_h�s��I@��Qs���i1sk�Y�Y&\��}���2 ��(�pRDl�܋�d��r@6E�)���7!d����r�S#x<N��.ܽJ����0٨���j�-8]mt�(�Th�Nbn������~���}vP��-����%�Y�%]�� ��tg#�ܥ�-���Q	.բi��>߫���Z�h�d� vW�y"nrʱ��g��x�ku���X��a��%��Ӄ���%�ЁXTV ƇP�U�Z���3��h��얃�����f5��	_�E�V�t2�P{�^�v)��X�?ȷ=�r
뫷[,@ Y�; �T���޴Gդ%��Ѐ�;qУ Z�+ܓ}4J6vP.;9LAS#.S%��[����ljA�j�y��q]D�)�k]U�������79����|`���J:��}n�r��.ט��[L��CĆc�Fu�;�+f���"��aX�^�� �+��̩ʻ�'�� �g�8�4f�y˶�t�?�c�|�.i��(r�
��d6Y�܂�]��S)!���[d��M����p�ʖN=K7�Y
�8W+�n��%yLz��:�ϝ�����I�(��Z�$= ��k����m�q����X�1��r��ͨ����,���q�?��ȓǜ	Ks�|� Y����8��\Ir���U��J�3$�YЬ��$����('^����o�(�K�I]����x9��-��-&�e�J��[�������J�))���Z�0�+P�}��.��f@-���Gg��"�^HdVk��Y�|X�f��$k� �i;�Mk��OGj �9��ǋ Ӌ�%|i�\�UW$�?Yt����aZ�>�4p̕x�f�asҜ+��|t|)M�[B�q���o�|�Sļ��T/2�j�\}*���`RO/J�f%1���͛@��;�8����*����Ý=��wg�u�s1����f��Aɢ�n���.�IO����@����e�i3�e�ZX�����,,����%�cҦ�<��Hhn�In�d9�6`�z#�؂%�'È�-�F�7��ʫ/:��@��q�)�8/Ib�-(��:�J��_�o����K�#�!�uJ/��A`��vvIj��S���%�+Uc~Evj��d��c��ꌵ��>�t��2�����`����<Q0����`j�{|l�����zba]�E��!�:=�νSdKy�o�/:,�Ald 9�돦ٸnG��;k�� ��l���P���t��$����y!r�KƐb�yi�5���ю"��	a0�p8�u�ԡ���p���T�0��#�'��
��<K1=9��/<MJ��/\��^ �����OYn��o�����"v���[����Y���ef�\�u�}�l�A12�i�.-�t�g#B,ފ�pOdn%�ؓ�"u?������k��a�1���B�*�+���ð���
au�Y��|��w�5Tu��T]f�}�Jº�- ��N��L���/Tz�њk�^���O�{�%e���p�S)BH;% �<ۭ`5�B�S ����Q������mx�^ǉ�����E�3���F5�*�C}r����bC"�Zs'lȁq�LC/['��?+�u�0���Xn�:?�u���զ�Y�S\N'���e�2�Yv���F��n><^}���O3�Z��]��	���+'}�G�5��{p3>�Z�&{g�Z���|���mJ��^/�p;5!�
%�}�g�`�"�7��HgkÃ�D��Zk=��Zh}��OO�˫NL|T�뿙���������8y��+��.����k����u��AK�ˮw���B�3�t�y&�����8n����ϛ�U�&�����ǢN:��%xN	�n�%Í �1VӬ\�� Q_9������U�O�m_NGӏ�[�vB��mJ�^��@Ң�K�X�1����!��O�B�S���"P4��Z�O�Vf��R��{���*����ߢф�
�==���F��&j��;7X���#3�S���UK����gS��%yf��$CѦ�7����������\ � �W����ޙ�������A���c��T��z���_�vK��]ݐ���:��n����Y�(���k����sJ�rͲ�����t��j*MJ\\��[����׸�^�.|��
��6xic�����p�#kp����][�V�H|�^��]qau��R�-��nUWO�P5o�#o�zm�.P���Y�Թgz�Ɏ�j�_a�Z1��׽����u@v�@��������H��ck��W.~;K+Y�/�l��3]jg�=�S$2�D�:��+�I'[����H��S1@�ѱ�k#�y���7A� �@kbN�6��:���ϫI�F(��{K�q�ڵ��)vI�6>�<�%�?�'=�cz��܌�p 1�<c����l�K����L�Abꑁc�'[w
��5q�D�)�E(U��像�[3p��|b&�~'�r�GQ�g�{O_4��ċ��f��P䰿IS��W��ȱ{M�Cʟ~D3K�0�)ּ{ȍ��,:�'���g�Y�rzR��ԇ�6┍8�A���z���:����mJ�&����Zʺ�B~۪���=L:<*I�z "0�"g���oO�~-ɥfw�csQ3�DhOʰ>��KGX�`��P���ZY��m>re�lÏgD4�7,����0oee�Z޹Mw�2�q�,N#4���6�3+�����O;���1(���)��~v�C�UL�Cj��gN>�ݾ��}w��)y^���QD��L��s����D�z��	�������rS|m�flC��_9�B]�+��Y���&���+r��&8��ϫ�}q�q��Ag��a��3�⛱Z(S�����r��p�9e�|M`�@;`�?����B�Dg�w.�A2�d�,'�J	�e�D*��wbT*45��z�`�C�{ WSRЉ1k�b�#��zN֨j�g�R�ȮR� X��=5�ed�;� �n�?:����=x+�AU�h���ˤ?���a6��7�*���!o�lv0�ۧ
0�)V{�xn����%���?�.xbtӛ� 
%.}sAN��k�!������p^^���Į��EYC���j���R�7Z<?��:���QK#3��-c���}Ѐ�rM%6ȑk�� 7M�����0HR�`(�[�"�#���-�Ε%5������YU�K<��n���,ֳ�|zp�\X�����6��jOj��R_�/$X� ����eA�D'//<���$��l�#��ݳ����C��A�C#D�������?�qD[�A�����xK��k��1�O�է�̲��Ջ�}އQ�e.Q:�HJ�Lx�|`������oT%{��C˴>����%���6�Ꞇ<eY/μK@����o�&ce������X��i�,	m��k��}^�h1s�K�n�>��М�I�]k>_�$���y��&Zp�;��#�v�o�+�����p��0�`�=B����������qH]RK]��_>O@]��Y�֦M�ȱEN�r<qi�:��Z i Q6��lX�%`;np(j�3�M�����/ii% ����il�Z��b9��8�f=�4hD�����<���:����Ma���!a��W��(�л��gV&NEs�ΏZg���Ż�|�˃�шj<�:�U��1I�aH�퟿,���Ԏ���"��N��w�?���\�h�y`��Lf#��m�*�Q�^��ngq8K4/��������t���;���
��X>Q��h��JZ@&�y@ܯ������ӆ@�H\\���%'6���5'������)�D$1����!�v����=�IH�D�h���҃����B��q�B;rQR�H��=c��EƤDdo�Hz�.Q����\�A��N�[{�¯i�۞�;��(���E��f}��vL�^� �0$���!�z$ �O!�Օʫ�T�,
�Y
C^��wۀ���O� ^�e�e��b��/���m���l�l��μQ�L�e��Ņ�ZS�ev��Zq=���nR���x���ݭ}�,����� '�R���CUPb�ã�X��5�ئ7���]�ρ��m#=0s���`�������������s) �o�K 2��}P���� &i:�����j�p��(�媆m��m�^���̃�O�b(OB!�3�qV�] ��.*�� :����G|n	����h�I{ɻkn(��5�mr��i�v�����W`��,��cR�>*�k�'G�ڀ{��w1�r�kʟB3�s=��*w����� d���������
�t�y;mh����d]��ٸ��������-Q�M�Q1WH	�A�x����;�#E,�eDD��5��z��rVX�������B��ܛ'�'����w��V���}*�:io#֕���Z�A&���c�LV������}������.;�/С��K�}�Tr�8�.��7��M�L��(����'�vC|��#}T%�J��9a��H�%��{忥Z�Ԉ�Ă���c��ּ�[����	�`�Õ��rb`�^�4m5���&:�^���������7?�76�%G�[�m���i\h����X/0�E�Ը��D���y̩�ܻ�J�3:�2#�> ��Y���Z���j;DW����7�q��-��N�'c]x 8
��a:X !�(K�{̀,U�K9|ZI�$��O���8)��"��0�o��po~���c>$���E�H�����-p��^w���~{A�#N����ö���󢉭&&q/�����<�Q��u����C6���*HM�:��T��]Zx�<�h>���1F��`)��T�ڋ�Y�o�^|�u�I��<��ܰ�D^d�@>����c!�ί����r���Y:��cʒ��{�˔�=D��X�������T�[}�R=�" ^���bV�Y��~Xm����RD�0G��O���ަ�9�� �i��ვ�@׉S�n<���N������҄���/�U�ИD�NiȌ�}d�Ɋ_|,��1UL��@tF;'.��_��涴��8(Vz֭׊8u�<ꨅ�댙�Xq<n��Z�[0�XX؜�c��<8��V�c���w�*�R�@���2���~" _�
l8 ���_�%h�c �Hu��K����LL��
x��L��9�>?G]�xϒ��^X�X�B��W[<yF��	��*���I�����pߡW��Q��i�@���#�h��3��~�8�����P�jP���1ſg���Ʀ�򫝾%V�G���$�-��sӬOM7�p�q�����jL��>��AY
��?��z��"H����(on��#�|'���c	3��bL|�4ڬ>?�5S�eQ4��UTT�A��~��l��w]�z��'��mʈ]#��!~p�L�a�,��+�س��kޒ����V&�ꟀGiL�*�{拈�a�?���F�l�c�2��敟J����[��>:<�iR�&�P��e����4���99����&�0��}����������t�º�����T�Uʆ�MK�${u�Ø��@`�1�{J��U�&Z��٧�-�V�.ϳ��~���A����LNJ���M�M�X�1W�V�x�����k�Ap�có"u~��u��@7�M�,������j� }������s���=�Ԣ�28�#f� ��������J�9x�@�ğ��P�[���\�3i��hqr�2��wx���l~l�*KV�{���c/��,��F_�4�\�ތ.0�,��U����8%��I6�^��U��>�|�G��r����S�l�N�x���Fh��|�1p�*��X^�s�Q񊕈�=����	����\b!c[�����{���XU��2��v[�65�Y,����z|M�у��������`��p]���p�=�\!v�7��<"�C��}�<��ܐ�v�X�:���s��;���4�33�z�Չ�_�B�����=8<�1�}����6@���Y��x� �D-K��3����ދ���˵��Q����"`������ƣ�!��LK�C���{"O�m�҇���j��	x]�~wI�F���O�|�wן]�|!����+v����$ro��5��/���]
yCr{`���Y�I��9�˳��W^����0���|��2�o9�	�����D�B���T���7��iK_�t#�Kt��1{n�-E�O�Au9h���,W7/y��'�/=�����;�֋fB��u�,Ά�v�8��0Jy�T��ޅx|������'�q���r�IM����������*��t����}C	��I�H��[�~?���3њ��Q�Y�'�<��� �v�:go��W+��V�¸�<[JyZϥ���_Y�H�m�|fq9�b�0]�9Cȗ@�rUk��wi��U��SPý�����'�蛥=�;�B�		��x(��}	)�W���u��]�F��Y�k4���V|fu�}|5�ה�y3�sk�B������ ����0>���Ծ�v"a�󷫼��.-����f�]�u�C�����?�tS�
_����[�Y/G&�Yq����cPa�TA2�Ǫ�����ڕ��?�|���jT���.p�0弛5�P���q�9�[o�N̟��(Έ����~����=��3^���ꭙ�.�АKb"�T���a��w�����Ņ%;�\�LYB��"L�i��L潧Z�o�2o��8��|�*�ǁ�����n{d��&����}VV"����*�"j���+�����>�$XZV��s�?�96>��ߗ�2Um��]�:�,�%����������z�����c�/"*����+�:��(�� ���w柽�����y�tu��%��������v�����
�X���tp�[�'����7������n��:�PO���}+������x����Ľ�2��>�ۖ�ou!c�v�����{�!|�������M6�q�������Tj�Ԥg�Gm�������j�އ������CBZB��������K����n�z������l�>g�Z�z�}�g7Hg.��ұi�ӐHd���م}���=c�ՋE~�),ȫ]�-�W�u�NN��u��"8�h
��y}@���G�������X����IXO��JSF \�8�o��Jr,���O����0��U(�@��y��^s�T.�s�n��/S1�Svھ,gsqÛ�y{6��� ;�r���������c������X3�9��s��'�p�1p����36:��9:�F~n�jd���*�qWo&��nWp��]��S�+3��L��	�=|��]�>�-��M��]o�~Y�U�\2��)G����"��`���d��=�`oc����+Wc��O`|�<o��U'�!�� ��c}a��\�(��,3�g+h=���ɨ�L�I�w���(�k2�A��(b�FEj"�&T݌����c���F�ᱣ�cC��+K��4#�� b0nK#65���Ǝ����z���Ȟ�0����o^5獽C#,�¶�bP?	�j�R6����Ց�s�ҟ��4ᒐ�D��CJ*Xo�k����%�<$��Ƹ��+��(O�s�j6$�U�F>��.A�\s{�7%��yy�(�)l�=�B�=���=���y{�e-AxrG0�Q�����k�*��a^�]��f{��砗�ܪ~H_j�l����lg%7��oʠN�����]��~�zywhs�*F7�:��wh�����d� �ϥp���Dk�5w�I���N��N��N`�\�n/�,�-V�P��6�42���&���o;�	�GY��t;�y8#K�8�	�a���.��&ێ�_��<�ir�׊]��;��\!3��z�l���ptG��)rI��֢A
�
~g��VBn�B�F:�L?�/93�$;�����dN���@ܿ'G�5��7c�=Mln��g�Gw��Ǽ�����M^����S���ɴ$�+i<.x�C��u{��:p6� BC]��LBFBY���pa����y{ȅԿM�]5����[Ն�M�������4�#g���X�U�fg-ߞjܞ�8[/�A��D�樉�$l�̐ۈ�m���r�~�����������6�nd�/u�z��߫Ȍ��6?�
A�['4��D'���e\�l�:`��܂�����Dl����|~p������D��[�l퀻rff]�ן
l-���s�`*�����uM���2��I'��$R	C`��d������֣7�_*`@�6GQ�e�!i4'_6��(d�֓96��;H���S��N.] $�	2'�@��4�18O�W�n��T�	0}XNB0_��@��]0�Id�n�`-�o0�`Q���+��J��U<<<��)H�Ŕ�uY[��fw�}��������R�Ep�D��).��}���,+)=D ��v>�b
m,�p�'kp&h�-�4�0G����S�hmW����>��]U�wb�eb�����K�Vפ���{��Z��ͼC^�H��"i�}�$�;t[Zc�u���<˨���ͣ�Tkzkw���'�{!D�-�ďS�ꪂ9��D{t����o�9�̊IΤ���[Xj��Nv�d����x�۷�]�ɷ�	L��K��GX߶�¢��r�M
��[@tM�,"�-��a۵?�!�R��Hd�yو�:WO��8[��0�/S���ъ�,�dE��T�*���YBrYllB�h�./o���Kt���ۣ�-���T9x���'~��i��:e�K,� `�0��0�tȞ7=��m�vo~����O��,쁙QUkc&�S��E��������=YHR�
���g�n�lgoP�w�[�@�ɲ�B�������Ê�%�(��6��=�k��jg�V�l��K����JY�H�{�pp���C���2�"m��a�?w>i�xq��D� �u�'UB���ձ�L)�|�W�Qgs+��+Ԛ�L7M�ə�yD��,��/-�fy��O�|��d5#[3h�D:��U������	��+m�@,(�ѫ�?q�O��y���E�30/ �������BWS�Kq�#�07fhfUQ[Aǟ빧��7Z=��Y~U����IԷgaA�x��w�9=���-��w���FD ·2��4��so����)B5�R����	�'�cӉk����3�<p-��|k�=_x#�Վ��7��Tٳ����j����o�ShT���@_$B���|�06&����Y���#���>	�t���0���n��>���O�6�Wa�0�-T<
�(��}gg�ӵ�C������H�%|��j�ɿW�P{���N��o�ה�<�;��u�}_�j�]]���{�:��l��ν���F�׮�ec>���mӢ�O"gy5K>�}�`�|L��	��0�s^q����^^K��LY����Zyj�]|�O�^�w��v1q��'k���y�Qo�v�s�n+K��МI� �DQugd�F�����"��oBh�9�M���UR;�j2.kԷ8E�;p#ր]�.T�j0��E ���}Y��'[�Q��P���A?�G%P���c!�{`�nwP��1�&���{t׈����)��E�/O^֏`�?&�>7M�ea�y���J?6\��[�e�2�,�H ��5�;]�����/_6�,��ڮ)J}���*'6��س���N>�����0%Lz4ʙW�O�ȵ�>��v��d�@?B"����4�|�uӏk���6�b�hw�$[@�y�}�g7M}v�,V�����tQNd��?�!�ct5�w'��ZX4�4On�45��ka���@�Z�#γü�á�~���Ey4҅a,Zn�xQ�6.WA��?��L�
�d�A$Ғhv�� �uO�3y��9���L����_��Ĳ��F����=��ҧg&-�03����K�ӎ��| +Jq)ۨ��
X�u����Ϟu�hV]���ă������1\�Wl��@�!v�)m���B�J) "vMu#Xq?����l�fFZT�;����)B�"�����)}$i!�!Ao �����7�l�R;�k6[ݠy�Y�8��VEV^z��i�����7�U�@L�ټ�� W��.p�:���p���J��K����]|�P
~��N;(x `�1�ۊ������6b�;;��S�Mr���N�p}b�%N	�M��	��	�&��b���78��n0��=�;i��"u.�����e� '�[lR�D�R�a�F�zr��9p�����ד��U?K����>��v�:,���B���{b@��m��,�?Z�\Sߑ52C���� �ʼAc�8�F8i{|�X�$�U��d�*Rx�\�cY�z˅�ADozcǼ~;{"j��Ʌ\�8s�����7�K_3�m�q�b ��syXOl��
��!t����`�����#ܚ�/:�~s�^�����6�������wM}�W���+�L�_ฟ�DK��I�ڝ�2�ǃ�nb�2��P�����嘆'�_8�~���*�G͆�FYȸr��Z���p׳ċ����٭��C�8�?�2D>ڷ��]i��V7�������U`*�Ɖ�b=�->X<c�ւ�ر����p%���ʷ�kPW��\���1v$)���wj���G�����yu��ـ\BЕS�(UM����b�Xzz�7Ooiؽ��!$_�n��@.�"�X�\x8|P�:^$H�Z�����w��� �;���
���\���R%CZ�`X��-�~��{eu1�F}�H/1��z&%G���uh�����b,ZF%�`�Ob<E�/�e=�J�����������Nͫ�;߂��ƞ��+�߃sUԽ��K��1e�v�����"A��D��L	���(�j*P�T���m��d��P�}r�YFY�#D��~\��)I�tFU��slF#�`��m�h�Hx�^�(ke_�"��g��o�WVĽ^.��0�"9��7� �-�H�Y���$�*â���{.(�M6��gv��2t_�3?'����DG@��ڸ�j���Ȕ�m���S�y�Y�O�շ1�D�ٸ�A\m�>�K=�� �/s�r�����/��j$ow��:���0��-
�,6�&I�+ �-ߦ��уԮ�? m
~�F'��� ��i�Di���Ĭk~�{�7��O��/� _��-��;��z)�fu�	����H;�9,��	�{����Y��.�����! +&�f#ؕ�����9�Z~�����2Hfd��_��L瞂�
k߀��(-�5��B����]ٗ^������$��n.���W����H�<�������?3/k?`	h�L�����Pey]�UN���N� ��vGO�c�p{��@^\gȻ���&�oU9ʮH>NIj���`"����j��΄��	kňj��ͲǼ�S��$� ��q���*T��oŶ�ZT�@e����S�蔄�cPh����vnET���J����9���VX�M��[�J/:�ՠ�J�w���!=���#*Z����ץ�.];Olf�7�!�l-�pC� Ġ\��C$���m��g�c���c�7K'ֺ��R=F)�PN����:}���O�,a�TvW�UN~�%�F�����{�p��:�My$�FI)f��p��w�-$!����ɧ}��̊�à���(���E�AF���N�ICc�3|��"-;4fC�G�a���s$�㺳�s3�|ͯxݶ�u[�A��܏���sւ��z�'��c�Ľ�]�d"�m�.�IRS��]����C���������^�.Wն�2)7�yp�L_c��A��_��ԇ���G��PB�?��پ�#��s�9�^���[͇U�6~�m�R'B	hJ|~0I��
{� 5�k�h���"��C�#拧'
>i~L�
��z�>ilM�?��+���I���h?�!���7S����R�6�'nK>4�IF/I�gݹfl%`:�f�T<�W��.�q�::r��"ϛ����PU~���P�W����9��3Ő���f7\U}��h&�x�S����N����v
�y��;�g^۠�,yl��`���ʸv�dK�s;�h���������K�Z�#_�=���I��|Ƅ�N�1�|uC�L�5��ҀH�@5"F�H��DZ�{���9��h��,V,�}]E�y:E��������7�y�'�WB������OZ2���˲3R��B�/o��W��|jǝ6�1��<Y5��.����m���P5Xt�����p/�{�d��TWs~[c3�I�"�lUM�����Y�B�99� �'�[������V:�q�`�\���08�A��Lr1 ���R��{���ueTٮd��a��w�Q�{�<�a�0�zq6�R���ն�=��֊��PM+,��&QE)A��L���][l7g^�4�O�qC�ダ���*�ߥ�������n�V��A���Ő��ެ/�5D|a�_����L��8�m��$�x�d;�yh�]W�t��r�<A;��ߺ�ʧ"M����p��&W�݊����_
 ���G����a2�f(��-�2�z��t�f�.�_���r�4p��u4�/$Fo`z�S�U@��B���U�&ig�y4 P�n�_�u�Qc�W=n/9�h;�6��Ah��X1Ga��M��]�����^�)��kWH�Rl23YI�]��_�)�q�A�-�3��n4W�	O����z'}ї���FV@�]�F��1�Ms+ �<�����y���E.�&s�{�b4���p����x�����n��ǰ��A���5��oY�@�O�/-[vP�tҧZEt~�-F�3�Yz���@����_݊֩���Nt8rK���s-92)j��.�������%���<4����j)7B�k�\w�o�y)EQ�S��o/b�4����fYT��k��E:�IY58\�����|Jn����`M�G�������2�(Mb�ț�G|���F0�ϳX)u��_���
��;�;:�oN��|N�R�6K����w�ܤ���=V ��s"#S���hm?�~�B�c���s-�M
�0X�A	Y�F�#�6�I�T^s~��N���$�}� ��e�Q�%
�߈���}
���0&]l��_��o�ѯ��1�* �1b�X��u%ō���90���?Rwf#)��S%ʔFbڡ'�Fm~�==fb�0��PMᯡ�'㷹��H��F�IE�탓|�fw�[�>X�[ۼK&��`�
Y������۵y���
SMq��v��eo]��=qPw�{��Ğ<>.��/
Rf�v��vms�����*�%ƥF|el0\_�X+��-��Z����:꥝�˸�E���f˾@�7�%ˬ������h
F�U�D��\��^����l�`Q�l���%u���lAۦ��F����}�>��~�;KL8������ oto�*}��-���@��A�vm��m���}玏���w���n�K��)	x/Pëg�u�q������hB�����b��w��*y�\�ٟ��)(3!չfSƄ�u:�j"�� h�?��W(x�|uz���w����C'�)B�``oݺWc��X���߳��<���������P�
���=��/_~���F�]�[�CiV[j/��u\�{��3X�bd��.cP�R3bM��V��K�6�l&�>W.�a���wj�1�ֲ�����LP���f�vt��{(���aHr(_��Z,�9'E؝j̀��і~k��t�+�89��*Z֙~� ��͌@��Xo0��E��X_�������D'ڼ9��c�
C���ˮ��M�ޫr� �C'y�M�1����i������f�	�����7&0��{p3�L�)5a�wu�g����3H	�!��?gҘ(�q`�R�ɇ�5�27|���)Z��P�bp�&4'�V����C�x�/�5��lX��gS�`W���Lz��
6��bQ �4�z�T�����@,��TLg����[�z�PD��%D�%f����ڵ瘀n0\+g��<c�l�������%�7�~N��A(351d���.���)Ӂl��DaA�/����Oy�2��1ƾ,i��2*�s�W.KW;%3x���0ơҽ���A�%�O���TdG6Xs��X�H�,,���ڂh���v+�!��l��e&�%X��~�_��� ������>�5���om����n�%4Ja�P���R##d�6�jG�"*�$��q��?�~F�a�=��wB��X����GK�(������j{��e+�:��xV$��i��R_���w�]2 ;�d����;d���\���[�]�u#.�m����>��ʇ�I�PQ���5{�[T���=i^�KٕP��W*@c�:���mU]6�}�ۮc�i!�W!��lB��C�3=������ǒ��O%�����m�vL�ؑlWG����7S��^����3����)|�Yh9�c��$���[�&P-�u;ݺ�7�R.��E9�@N�� ��L̃3ϧKU�:�����3���N�a5�'�"(�e����OL�����H:>Ó~��[[��f�Uٷ��7��H�Ѐ�G�<���▙�Q6u����p��2�'u8��1�;�����f��e;��p٧$7�hv(ӈ�X��^1��?��:-,��"*U���Y�u�ܐ���fm�Et���}@�T�U	��|*~Y�A$,s����lGf��t�j�u�~��\I���Kt��-En�:�'��\�����c����m��J��ã���wM�u>�]�2(J���䜷��4)�u?���EZW3�]���W������_t���eQT����������}���c��ټ�uؾ×w?��#��j��;<\��({����l|]�����/��a�*w�^�ႇW`�H{�1�4_��0 b	�?V���I��#O�u���}��F7��^ui�����
8�T������hIy��Ke�mQt�_/P1���Q�;���j���K����}�n��X cCㄮ;�(��)D��cSr���%r�)�	S��S*Q�mMd<�����׹q8���q�r�6xx�]��z�A�����7���8
Z�������[k(��_��W�k~b�f��+�,>�2�hWU��_h������E'u���Ht��u�2����7n����y�Hf����Hbݶ_#�F0�o~�}��i'���~`Ct@[�Y<R}���o��u�����2��	o��䩔���+�qjޮ���X��๶9CjLk�3v$��L�s���fWYy��<M�oT��n�I�6V���m�nş�	qMvS(��g{.P�/��Q���?��#�%zN�K�����!y=K��q>��1�<���}:}QR��X����ѷ�����I`b�_�"h�"MW�JX�8#fd&�o[�M'L�bR>��EQr��w�B�,��r3ʁ��ugv��^�)��:�b|ڗ�Z��'�@�1t#;aF���ê`^��P�D�����8�l�2�]HqWa�ňQ��h*�� Wzm<��<yd�
���S9XKɕ^P � ������C�Q�����`4[0 e�o�hj�n9R������v�Q�"���8��}�auT=;wd�_@GM~��W�3���^����<�}G�%�מ��YO;V)Nj� �����AqPڥ��^�%��9�3.)3`MH�������A�r_(Ťy��-c����������K��bN��� ��� �Ή�XG����g�垉��=IJ�:�D��r�� #���1����<<�������2 B��_D�9y��+x��CG�9���X���͝ɲ�<���_���ۻ�C>sb�P�9�bp��j�'f��Q����Ic^�z�����{0��Χ8�fU��҄7ߧُ^.�~p��\=�~�3�O)t|$��FMDfV�!yn�M_��P��C�'���w�x���u�k����(ll:�@^o�z���O��6Ul���)�g��W׺d��h@\�"�@��@d�{F�\�~�h�z�`��(8����@n�~�Q���M����G�q�\�JBr���C���~*�?+�� �uW��g~p�&�sh��_Z,�`������K�W�h��C�՜�|��;��ěg܁+��jQEU��r�Y������^j�<>�2���݈��~h
I�V&� "SRE�g�%��Gm���a���Q~�0���+�!�����K� y艡�$�YG3�P�{��>tdGSC�p�;)7�;iGE������5{50�@��7��hG�_����{���!������1W��w���>�|н�&RWJd	eJM���d�?��K T9'Ņ���-�O�*x� <�-ҽ�+"��s�A.q{��r�{M�-P�	�O�y0�I�u���i�=IL�}v򢎲���	���Ɨ/�P�!�@!�?[�M㹙l#}>�`U�~�$�Lqw�G�IS��] �Spg)���A�c۴��p�@$xB�����ht1U��:@�����#�*����g��y���k�DB�+�l�kx
C�T>cqܰ�Sd��:�eB�v�i���Ƙ���O�ȟM����3��ڷ�!���J�q-&[�[��Г9��TE���i��* ���D�{T���ն#�ҕ[�@<���n�*�8��s�m�����B�2�pD�S��C�lf��a9�,�P}���C�0(E��:��ˌ���C���5��Fe����&�_z�R�e#�%�I�ք*�v�+$�S�7e��ۘgs�[lvsD�i\��6���{OO���5�\!@�Q�T-��<�7-*��n�<<���Ud�g�����)̀�V�,�P��|{>�I�f)�(��ϟK;������B��<}�1<�9���D<|�0�ؔ�'�&�1��0^(��?��.Q3��˩ӂx��=zh�2���4?&��aL��P�?�PQ��o��`�l�L���D�A �[�=D ,K�,��Ds���>@�ޣ�`R�����8Ƚ���t�=;����\�R 	�"�F���EA����<�zLY��G!#a\��
O���j�=�Ӻ~���k��~�ШΘ[a���z�OU-�jY�;${y�ѥ��1--��'_��X2)>9),�k�%�f��毷����]X�𱤫\��y�x!z��l��
��b&�y�e���L8�l�Z4f���3�D�M� �E�҉��Y(�\"ͳOz��#��ۄxԻ�����Ӵ��C���,M���<UX5�%O�ڈ�lo��UU��%
T���7��������_�y�yPZ��$����o&�WvN�%�Q/�`��O
�����U����x�S}0�so�&8 n�R؛G��mz�oOSyND�7�|�a�4ko��`�����)R�ǰIˑH3=�p����R�����ת�xmm��� -Y����� P��>`�0q��0ڒ��xo;�V���զ;�i'Pg����ÈG���[1Fw��b������%���/��!O�q�*�o���u�
��+�$�F��tH�گ 1��X������?_T�'��`eR(�ebSq�g�Z�nF�y%邾�����C&x���kU�����ܣHM���9B���i��*.�*K��s�dЖ�\q�ڍL��W�����xa�w����L�����̯��R����N��������5��s�I�X!t��fU��2@�Cm��sN�џ��X��x�*KO�3� ��Vi9N��� X��BOa!>j|c"�}&��if����5b�C6��j�ɑ���=%q1#6�˲�Ȉ�S2M5��H��8���	��?�AD���u���'�,t�&��`Y����}�:���R �W������q�<�eeG���R3�����l:���$��$ٟJ0`'�����	&�0=�ⳋ4{�@�d����&�u���.�-�/Gz��K#.�rh��",��'��Roa��?�0`+x�@�w��&��r����;D�h7�Ę�����{�I�����k��Vb����%�ט[M��7$�k7\�����A�	h ��D��F��.b�#�gu@��Gx�<PC{>uxK\�-ፎ�*�k���;އ���]+0��^��8��,�`;X�qi\��/�Q�̶
aRa�X����㍆47�Ym*��H�KW,O�zY��4�˜�H��^g���A��<��)�����J*�Vs�}:t�т὘��e���L1I�D�1y>ܤGK�V���ϩ�2�OCP��2��y��h4�1��J	qīCf��D�Fv���`�a��	pX�} �U�q!�����LZB"�$�f��?��<�8k-9���S��9GҪ�Ԝ7̠��C��p��.���6Г������=�>�p��RQ��7�g�e�:?���|"w2��h&m<3`z�q���:�B��(��c|�w�Qu~R���F�7�L�[6�C�`���<~�0f�W�#h�iy��%<2�9��L-6�u��F�pa�h����M�] ֪������i��T� �z�� ���B�coV��Z���[U�k\ub��/�HrA�ӡ){QSt��ZfP<����T��1�{�����`�/5K�<�G��"�]����,��s�c8�'�\N�pRu-�x�6�����Cc�O(�e��/ŏ8��ZD��V_ߑUD�2��E���".���$N�A�t�j�)Y �_���՝/�&�+����S	٢����g�TE`Hv's�w�c��@���K.� �M�9�Z�T	�(��g�Re������!����6
�?+'g\�d�G�par�y��T�Uz���ɚ\�T��l�Hh�h�}0�쥝��ěol��+�v}�-��rz��6={顗ƈ�+���R���!����+��}u"+�Z4�<+SV���ό��7��eI��߮hg5{ϞJ���	ZҰ�跪Ȥ�� �ݡ7����;�-��?+jɌ;�������	'\8�Y�����5%��7o�.t�~2Mp�a��mB������nd
�F����c		\|]�y�jn��&}(�6�~���O�9�H ,����5V	b/q����$��9Č'���(9�E-�;3�+n¢J4��2�q[���&�#�YˌS�/_*��Y�aø�s�����i�[rF5�[[9L����@<�y��VZ6Z(P�M|)��L��*g7�2�2�WD��̐���8����Y���#����+��M.|��+�Ay���;����X�faE�o'^=�S��(�$�Z����B���>Ξ9��v����Ih����f�w�rS�3��[�2��` UUǢ>��GB\�m�zx����L�7l@f9��"M��_=�
hv�1Lr[��6  xt���7C��^݈�\b� E�Aj�4��ʨsy����.�S�z�8��oZ��Q����������#O����a}��~�o!����׺5$��Gb�K�����hk!���]�������� I���:��H�W�B��K^����>�eO����?�DKI��y�?I�m��x��� g�@'}I�	l����闁�H{�9�[^�<��V�5�c�C�T�����5/�Xi�3c�WU>�~��u�����[�����IE��I73��ZS�G�w/�+�i�y��u�p�"�E�N56�2��#�}�4 ��-�J��Ɵ~	{;��^>��X�?@��!_���|��@��B4�w�-�'�cm���B���+��HI��wD5:�.��
���7I�!Ϊ!N�Xԫ3�t��Xf�͖}�d��Xz��KHX��|Oˬ�� ��D	AHz������t?θ�ߣ�>h�\��A��<a'C(<A:ݏ����'	��	aj=���Q�N�~y�|`��'�-ޢ	��5�^���6�@���&U�ϕ]��JG�O<ѶwV��L�$8�����Q�ڂ������`g� '}	����̃krI}yH���i�Q�C�g\��27؏;ռ,�{oY �P/�������$���Q��1O�M*�*fi��7I_���Š�1(� g���-�!�;��ǻ7K���~��6�������|�c����m��B�� '
�~n��X��O����w��H��;�9 �'+�=>�y�+�'�d��0��`\�U�3���>v��#�õ�|��3f&��~��	�6��t����(����rT]Y����Q���O�ʁ1p�Z,�r8��t?ٸ��*A�D�G��/���S��!N��W��y����Z�����|̝���,i�x��W�a��h2��4=��߿?��ś���`0!����]�9;!�-���iC�J,M�MY�}����a�gk20C�������:���: �RvFH��:��eD�*�|��N�zV�dpP�I�,(�P�xKs�Sf%y�?I��-0=�"�!��4U�=u��w闥�ܣ��/���:;��	�Q�� ƫ!���U�V���e�Ɵ
��O󉦸��:��j�AS/(-���rJd�ui�c��>��Ԣ�IK�4;��	�;��j�zu�y���Nh���<�^��s�>] �������Yޞ6��V��D,{�$�"5
4@�~���p-�z(2�G�A�6�E^7re#
���)�ِ�6̹K1�O-�Hƫ94橇�����3{Z�@��޹@{⌵��]��.�2.��p>aҐ����aO��;��~�������̨6�~L��^2�*	�I��c DB#��Nb��^��(�j�\n�5Э�,�0n�S�qw����y5dǸ�/��GP'�W�&r��k��Լ�ϪE`/Aq�0 �_�'��c�Gu��:����'��%����r������8�u�br@���ׄ��@|/k��ƗRs�����)�;N!ۃ�x<��Q/_[�7��FB�@`�!W4������Mdm�Z���5���į��Җ��7�7Y(�99�(�= ҇���)3}�����y�vˑ��:��mN�觎����QT4��N;0�p�K�e�8-�m�Wf$�"�
�Z�K]E��/)Q������鰢I�_������P�W6��*%G�����Z0�������C��~����I��X��x3��tC���^�QCN�Eu^�_q���6�{��U"�2mxW-��og��p��750������ux	����O������Lwqeh�	��NT(����|���Y%��!��1&Ǫ����rp�t��m�=��/:&�\QXvg�AC�/��;����|��':�4�#�IT�i�J���w�0���f�N2>_��h1v�]�J¶�n�9M���{+	�[�#I/��c��X��a�4��$���c� [-�N�*������)B�Vf��Wn��aAg����֩O5. Eq��J.5��O����,'8�f��A)'ZX��U�	��
uƁX�F}�>�]��R�s��2w�7`�5�������/��>�ͣm4G7N	��$��x����w�`�e-��ܮ��<V2>��8]���f�vx���p��x��'ֶ�x�Ś�8���Q�9��w���i`>��iqH�/.���p8[�jVE1"�L����.�
U�(�O�B��u�����8��=�2][gb�����Xژ!?W�^jv~̰�;v�ŏ^�z9�''��-�sb2�[�;�VT��C�Ҙ���Bƚ��yq�MXU�u�����|(���ok�������y}b�Uv�׋�r�%�v�(_��eη�4�Ӷ��C��^4𕓬7\�D���r<r�,�p��Y<&��A�VS��V���]ay��wV�k۠��SI�?�l��3��	�5^��Z"����U^%��k4�/���q����q �}a}���%�ւ�߇�E�����ռ��c��v�S�M��|ׯ���9�`z�$2ѱs��|JJ�@0���K�H8�����|��#����x�OGó߮�G���4I���{��K�gX�?��~�1�_NmA��2�d�����c<�,-�x�7Qŀh/�}����u�A�y���)�K(���U0�V�#g�۪�ͧ�"�4�Gٯ`�����T��$+;��Z`S�Pw���		ko����Ys�<L��%X��ڗ� ����H�8ןA�
�/-���6�����oD@n�������7d�Lْ�ZJ��g�8� 6o%��ퟫ��fDq@2�KD�u�Q�]!0Fqz��x�Y �͓��f��I<|lw������_=��r���d��X�%�ق�r�Y�T�"<!�2���4�Q���������5�6�?�$�z�Ď\�ٮ, ����=������ ��T��u���5Ӥ���8`�fz���|�n���������7뀦��T�Ƥ��.�
��xsi���e���XB,�{R�t��5�o[���t�%h������I�cf��Fw���J��۲1P)�>�Y�X���Y�+� �.��m8��.��k$ߵ�����}�L�)�\��}{�����Qs�����J�(���I��׼��-��Пv�Ҫ��vPP8��Bv�`�Q��j^�!9P>B�6h�B )���%6gI��Ff8n����	�Ň�rii�����s���C�}�{��m\���K��+m��.�SB��L�ڵ�[��D����n��X6l���9��nO'����J�q1��\��F��CIy|~����)���4f��*衂�[��2��r�~u�|������;�ujy����Ǵ읕���/XDD����;U�+��_��n$�S���vv���T�����X"�O��鈬o�74�E_�V3����x66D�`���N�*��e�J���+1³7�dFe�O�K���Z��H��/�Ff��6��"�
j��\�*�bI �l>���o&����w��L�b��6�z>9�����00�#^�Kdґ��n_�:�ec�����ʲ��!�T���w��Q���]R��b����e?;�m�I(�������H��)�ikU�\�<)����t6x��l^T����0�u� 2B�G�_\�u�w	E�v�FD&�"�
Ƚ�H�V~�:�h<|�7���Bg�}S�L%fe��ܤ�L�p�_:�=#��J�x�&����ZL�ߌ'���B����W� E� 3*�ﭥz�M֛XQq� D
�7�r��0E�q����UJ����Z��<;OG!F��cVY��B&��f�n,N�B�ϣ��׳.��;����澸�7Y��v;�������O
M�L�^��)[e��1$����1�ra�G�i��*�])��Ns�2���e9:���C\�����ԅ=�+G2"w9r��F yUQ����p������?8�O�Hi؞�z*�_�b��&7���R~4�9O
(�_�� �L�!�6*�h�����h�g����?�ڶ J]�f����g�LO��v��{Si��@��OU����60DI�~H��\���I�u��^c�.�XM�L�$�qm��5w|�[m�6ak׸�R�}1����_Q{��������͌��2[y��-��J���&��f%[��b�N��7��R�N&I�.xH.E5� �����~�E�c�"*�ϩ����udcB�%B�U���Z�?�Z��5�Tj��4Ns8퉹��U�m(Qy�5,:��]��\lp���p�,gC0�amo�y��[ϰq�p��
/)g+􇙔��"�J֪%�gs�K��fKU�"���K�}�#�I������u�D]J��V�e���?�D�(�W9M�Q���Jq݄��vי	������\;��3>�Ə�
�w���U�G(��u���C����ׇ�V�r��(�e������0�3�B��AeU�|�g
E'��OL��_��F���=i\�ĝ$�[�hC�u�hM��KY�ڕui����J�Tie���V{�
�u)Bu%B�"�6~�U�:��r�|���}f��y�����m��Kk
�գ��B�~۾Գ!�fdk��4=��v"����9{�+��by�F}�l��x���C��.(��ܸ�
O�1ݚ������w�g�`�?+��Ƅ�����>�����bUb��!� ���QJ���[�q�Kb��[u��Vp#c�;z������+���W�����ͬ�S��_�±�"M�C��o������*0�sw� ���j�v�-����>yMg�n$��|⃸ti��S*i\��/���`��ڵ�=�����g�d1��]�˝��xU��&�MG��|�d�>�+}�ǃ���b�ya��̴5��%�˟�FR�n;E�#�v�3}��ݚJ��Lc5?��V�@�xP`����-<� �`WQ�x�S��xw�M��sA�FV��&�x;C �*�*�V׳9���p/\)��ƨ�)��#;���q�x��v��z�K�u�8�����I�u�׌����d$����z}�i��+{�ǁ��R{E~�F�5�@,�N4��i_�ǫ�о"�u|WR�dM�`�I���`$)�B�Ճ��t�\�^p�3y"+H�9τ��4�n�E���C������Upm�ѠQ��U����ifru$-���f�Y9o�g�,OKa��`����-��L[i�c���B�=�a����3�{6� ��p����+�r??,��=wh�z�c���L�Gf+u������A����zKP�C���A��Q��!��x��f�qX�5K�<���/o�0���85#�ԝ� �����S۞����8ɚ��u�-q��1h1Y����+$�c���V����^�d�E��Ñ�.�PI�!q�gԥ^����'�V'���#m*��NWC^��[��!��#F̙�;�w�$��mf@>�����y(���H�Q�U��*���Y�*�YԮ'L�t_q�yЯ^�,�Ɖ(��/�F���P��Q��3�m�䮹�o�}K

��*�uQ��2���+L��WN�A����0e���1�٬Z��"�cZ�n
J��g�R
�����F��B�����o�����\�XM��α�e�X;/��c��@���O8�ic��P���(�B��+;�ʗ�]7�T�u@*"oG��������s�\R^���̲-�8.��-L�GeT���R
�ˋ9Vs������Ŀ���:�d!�kJ�u��q�E0���.[�Y/��^/}��󮘾�R�ܓ��P�V�~u�?ö4��5A*���Ɍ�����<��Uhj�Y�;���*���)�c�X��1�U�����Z1g7�p��#�1��U:�C%�N��5�(�cȵ��񦰈?�ӭ�w�����������䵔.��p�h<��"(/u�(}��
G�g��T�[�I��H_��7�A��WlK���O��,*Vh_�Pih3}�7_�LM�t�hZĽo��)�-gI`��?O��W�Xf������^V���B����S��j�y,<5}�W ����'�Z��+�ψ@]KK��Ci�ۑZњM��/��*L�r�>���M S3�G����	����`d
��P�O�$��L� ���4�Ó�3�I@�.Α-S�2���i艶ͥ���F�T^Y�MtOL�+T#~�	�W�����!�P�;_�7��~���]��X���5p�"�>"��<�+����i �L_ظ�Bݬ2�v��ٳ�[�ޅ$�-��̬7���5X�~$�s�ʓ�C�����y���A�Fn�e��2����,JI6���.�
�t�Ø_�����0�5Zd��θ�����`����<�X�<�
PN�i�p_?�WK��~x��?�qO��7�P� �������oV��'��=�Ӯ��_����gDY��%�|��#��c� :sv�5���0�e7��F�%�|��kZ�)ʘ\�j}I;z��RvM� �eQi9�==�Ǌ�Zym�ˊ��g1gq�y@�3��c��t#�Ky� ��oٗ=0Mq�w�MY���ݩ��L9�"D�m�>3����[�~�8�,�M���^��Be=�	��'�~�8��F�D����}U��G�_�0>�(CJ�j�{�Ǯ��$��H�_)�V|����yo�,���ԩ�0fT��`J��w�	w�¹��u� ]:Q�뙏�ޛ�0�w��X�����|��k��	��%m�@��)�W��rnU�ӷ��¸��m��]���ev�8/��2��«ǰ����S�pK�
�q����f��>����%H!-G!�����/>��ok�M�xt�՝_�~K$j=(�PK   �p1Y�N��i/  d/  /   images/3825b8ca-e3cf-45cf-b79a-668c63877d2d.pngd/�ЉPNG

   IHDR   d   �   �{L   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  .�IDATx��]�Se���}���ޝE��+b;zꉽc�J�`�,�)��,�z�X�� ���g��*uK��'��?�KȆ��K6�d���d7�׾��i�������O�n*�R7�L�F��&��4��4�I�MG�1J<�Z0H&���h�LV+i���Chi=�`�9���Iުr��sW������(f1�ɘn�!�t���ǝB�O����"?/#����p�>��d���c1
�m���i��~������\�~����ߑ-N�-N�1�%&�E�.|�?��g� jgI%�K˨욉�t�D*9�J��|yN;�b�M̤x$m2�-����=��wY��XdY0N:�A_�#�ټ'�1gy�ZZ1%s�D"�D-������g�n5P8��w\0�B���%fLW!�0�g1����C��}DQ5�SX`F]�j��#I'S����A�XD���~�=�n\|e�f��W���vr�qh����/���7���	��;29��χO��ڕ��X�cU@d��*���\I&��)��83�IK��q�r����f�1�GK$*��~灴�G_R�j�s�1�gf��]BU�<F�vI�U���}��Sݥg�l��L��0e!3�X��r>���K����>|�c����'c�ۯy��D@J��ke���P����+f���?䴯c��?�@p^��+L��✭��@�`HVI��FȲ� �f��YE��C�\E�m�K{���'U�9�֝1��Y���	z��I�j��(m@k�X��� ���៯��N��ɫ��ҡ��)�q5=p�����7��P֔Kt�Wƍ`�CIC�<nce��uX5�"^�wqN#���5�Y:b�n?���D��_��g�Tz�����fTr�y��z^�fD��|LS��gF�O���";���+��c4SI����d&sY9��N���*F@O�C�����g��b�����N��I����N'_�L{?�Y�Sp��ύ�*펔ƫö����@�5z)���Tz��d�rC��<�Pj��]��4˃gI��8�����2"��8ct#���"5�>������=ؒ��c�~d./'�|ҝ@��N��=j��R���-?�?��C�`�`'�d�՗,����W��ˊ!X������c��ךEٮ\�AGR����ǜDČ��ly���3�
^������7����FɇY���}�|���\cV�(�n��c�7`F���"�,!��voۢb���0K�������03�	�(������5��Bp���u���?)8�MVY� ��x�p��z���	���Bg�J<r	�-�a�2A.i6�9e|.~���"�-�����9�V�����.�3�>���.K�^��E�)�*~9��tF6̈�z��#�8��`аEU��>z��F��Qx�uѫ�_VH88�>���`MA�Cg�[��}���Gylp�5f�b���x�d��&�.��ǡ�R�īDYCA$�#ψQZ8_9Pe@��?t���Hb
[j0������KZ�!��/R2�2�I�����'�������?k�>��/	T�Z'� ����^%���d��w��_�?�6\��_�����Y���t��GR��w�w�X�`P�g�>Xo��P����<c�2�����PՄ������/�g</�|-� ĦI�$3�	+��wS�Y��Q�l)�7������+�b�=��~"Y�j���$�#��ifܴ���
��ZX%���ci�!�%�b�4=x��?ɟD����"6�p<��M��:,���w��a�j���Qj��BQ�ĺP���=��׭)!�9O�ta!0B'�������ﰦʒ��6,Ϭ=6?d�=�����C�
�8�ܗ�����.�F���t
bS�4r�;R)I�,��e,�K+����!��#��
P�x[��-��:�3�,��d'���iX1_K{�"|�&�?5��2��VX2;�s1��%џ�R$_C�UW�LrD��!F0a��J?���[J*P�O*�l<v��Yw�ۣ�a���[={0 �� V��4�|^
"B���\�$_�e�� �29�	3����՞SL����zrMV����(��"V���]C��O?���VGL���/��ˀ�]C����\B7^&�>��ƿNV�Eܜb�����k2�e��@-O?,�i��Wr{
ߟK�9���kL�K�r�$VOӆ>���RUM��P��Oee�̢���Ч������)��+L8� ��:���{,�O�:�8�x� .ͣ|��!�N!z��R,ɦG��w_����:`k%�r���
n��1�<�,�V�/�q�w���#}�X%)�����/��g
�UL�J�7_L�ң��-�w�)��Ƅ��yAWzLX�lfD���Le�Ä�a��ЉA��? }�4�SR�1�2	,�`T?�"���	r?A��;�Z
~��YG����b/#Ø��}LX�2�<�98D�E��}C��K���eJ
3�ӯ�1��\#̬Ki���o�~"ޞET���}z�d�+�(&�R�f��M�:`&byPGK�x ��K|c�QC`>��������"e�{ ѣ��9�\Ir�?	�V��yrrp#aꔢ~M��QVඝ� 	�]�Rpp�`U5)��
�#}���.�!�r��@*As�*I����E��m��S��J�	�2K`�
��9-&܊xfA\ż����.�Z�(�� ��1٤�`��4�灇,�xf:#��a��T�J��/K�����v{����Q"�c�p��Ą����y-�%?�հRJ�	'������/M��[��s(�;���{�fJ�(�p84��q�*Q��lQY�@�o����U�{�9����l�����K3����61a�f�ɼ��&��l��a���>�q]ǜD�wߢ�ge���L��TD���������]�Zp3�^L.Y%�R��sL�����fN��������O��+n�t~����w�$������+�	����,�n��}�h*9�"����z=�<��Xl�S�&����ܭw����`;��9�A#/�]EX����\�'�QǓc�}
.�C�ET�N>0�\`��@lǺ���2�1��xA�$� fd�ŸiH�!���G�_�Ď�۬�g��ꩲy��;�	�;�Ey�]|�,u�nU$އ-��sN��K�����e��S�&��"���]�����(�!VDG�7L=L�u%����@�R+���z7�:��wD�0h�׹U�g�D#~/�V^,��Dt���|�L����ú2��VasfVVR,w��^:`;��EjoH`Dߕ˩�vuN����nџ,�k�B����Px������I)1J�Q胘�w�5RSa�)`FC̱(��;��<�8��ҧE٪�.~�z��o�Ll �����������w����1u���o�]LD0"��,*��V	]7?�@ǖJ((ް�c�"��\�M�H�_V�M��+� �.wf��=�R^)%������+UL�����(q���ԱdYDYz��q�0�y�R,j ������t�e�=C�Pb�~ r�:_�h�U���D.&Q���$�z�XCYz�t��1u�86�h�]9����L���d��RKaD��P��)!bS�\���sO����m�]Y�Zڵ�c,�,�ȆXD'I%�bK�@�+T��&��;��V'�����{� ����Q ��%cx@����
-m;���K����.�m>z�"����ot@l���6 �,	�
I�*qQ�)N/[Y�u�����֩g��;�`�b�y��d���PJ/��\G��EW,�v��kX��Y�Ml��x��� 1��]Q�v���[!\�Hʏ�C��2WTʟ�/<E&؜֩���yPi6�:�`Y��s�^xZ��`�T?���25N�q��Ajf��RSM/j�M�JV��~�W�PNH�Cji�ɇ�}����EV�gs�}�����d��7�����<^҈�$�Ҭ�H�(u~IJƾX,I%g^�3t�O�EeV�=�EH4��:��9��d[}���
yz5Ն�
����F/���'�����Use�����yV�WJp�|�g��A�W�&���6�N��Pn+��X��W��1�\�0�J
��}�c�hTSRJ��v��7_J	[������(�l����/�Q��/%��.uxXRj�ǟ<���3�@d�]M��������Vf%��&��Y��:f0{�(��~�=׭���ؚխ<[C���ҘիV��=$�wkCy;|͢�sB�լ�K/KZS#��*	�~���2O
S��n�<nÊ�vr�Ee�^G�cO��G�Ʃ��o�ă_�P�F+���8����-�zK�ɺS�$�	�St�J�"ض�Ar}c6sc�:��u�r>@:���;�;���ձQ{ۢ�[Yh%�Ć�g�v"V���V�bAc����y��V��}���fPd�R��Y�?)̐�;n��n#װ���g)�ޜ�N,\L]Y�����]�, O��6
�>�i� 3Y'�IiZ?����{l����TaЮ\��)��q�+����n��H��YE��?�P,���hBPx⺢�����'��9���>�JCzui�k�T�~�L���)LL41�p֌xϬs��=�⦻��Eo�7K9���؏�A*ｕ*�|�Z�{R�rzN���ƽ��@�bҽ�M;<���@�!�AG�}���Bj��b�Ah������!�S��Lĺ�@i�'�Ѐ���t��J/�N������k���)�N��]�.��sY�?F��}D��, Y���Y�,_&�*j��v�j�*(L�z$UL�*�t@(�j��<����Y�!�y�e��_����0�THXst$UO{N�碙3���]ry�?09���J��@YQ@��ĝY5�Au�t��b��t�����vx	(n�kY6�O�w����������J���v$��;�R~��2x��}D�p����Z���Rf���J@�$�� � ##~f�(8��%֞p�0�r�QY���KJڂ3��b���/�ՠv�ձ�k�yW�֮��\��B��%�x�-���|���<	b��ܗ\�Mecng�C�] ��C����A36a*Z���r�F\�
_m���֩��,�`���|9�[�C	�/ѧ/�X�F~��֎<H�-�IgJ;A(u�t�@U2ҫ��E�$]{���#�<5�W�D*9�"�?t�c��|�����!1��� lO�B�~�X�:%z�޽��c&���1��n�,-�|�Q��7ma^02:�� :'�YIK
��C��g�HB/D(������u���Z&�D�T|/<��֢�a�yo��E�Ϙ���g�i�3����;V����R3t�b���~[�<:h�V�����iIok.���O�ґ�z]����	&]l@�KSN����7,�UN]C-�Q��,[�r��X}Qe���O�W�#�]�^~�ё�'�@yycꈴ�FK<�NP�e5?|/��y�X���&3	����ؑ8j���F���zu0&�K%ّ��&����t�L:���E������d�Bl�������������;�0=�XX�E�}�Ѥ��E�Wem��}�/V
�R:�Rj��Y��`� �d��+�Uh%�,F�HA�"��k/��x��"��%���B<���G��~'M�"�lFu#�ˀ�����WZ�<�w��%-�V�$�'
������b�4�A���1�EV]��Bx���3���4V`Y)��X�����y��{���֭���Y�W^̸�J����^h�lq�$7
�B'��4��A���s.��������ϩc# �@#އ��u���{��Tu��b@�j�{"��(pL]��Bc��V��3�0=Q�	H�� �)X7�#�#��W�x��2p�~H=#���=eFGW�$�n{�&7\�JѲ���gp�7T6���\��Q@�̘��ԑ�PQ%3�	P�(�����y2L`�}��IMx����:z#��zX/�(Sj7pmL ��/S��k�m�����aea����Q�x�x�`"`
���-pL�,����d7+����g����@l��0$��}�񾗦K��c��F�l���UI��n�MT�I.z/;���+���s)8�M�����+��&�ԡ���L�d�[��L��� /+�=H�SZ)ăYv��T1�n��B��*����n�6��������ʱ��C|�/�Z�`2��N�-`ac��5�ٵ�H�m��`_��/��>4@��Y��7�p��G�I-��`�-��XY����\Dg�ۯ$&fc�%���te�d!����L=%%C`i�?��>����)��Z/9��PL��Ӿ�Z@eM���	��g+pj��nJ�P�. �wE�#��L�Y3Ux%���k껩	��h�Y�5C:JR��o��Ә:��dR����������cXJ�I+�Phj��8�?��'*ؘR�����M�qw���ƌ|��OҜ9�ݕw�I�y�~����S8� [k�	c�
�.o+�:���x��S6��b���,���&(�('R�SH��J}v݃~~c�L�a �4������(��Č�=�y������"���R��+��4�rJ�K��wx��s�^��e�)p��@j����U�>M*�H2���k�=`�O��`�Z
&�Yo~�$6Q�I�G�]�&�t�"�9�M��&+L=�J���"���RW6w�R�Fk�X#�"|��ǋ%����P(D�:��[6�!�{��޴+���C�^o��y1~� �U�LG�����sB�L6[�ٺ����(���*a~�Ɩ�F4��6�i��1��gv8L�K�'+�VfJ�7K�ke���Ri��z	�n�G�a�ѥeaa!C2�Zר)<�'��y}o��qR��b�U��z�|Y�3�ܳl1�x �|�W�"Ӭ��w"{8���rf/QS"��$�"����7GS'yX��{ƚ�JA���Gf8��$�VV6��IE�)N|��j���y��OJ�!�&lv��a���)
��0��ׇT����~!�*��7Ty˽�=�����AK��V�N�T����p����<:�"6�0<��>����m�U�)�_��.♌�H����:�� yH�@f�����@Ot@@"d1����`>�[$��1�`i1��/э��14
S�iR�6(�.�Q��������=�P���Wl�z</k�Ҵ����)���m��E��`#���5JE���$Y�� Kt���U�a��m�������$1"I��TC�4�-��Z�4�@**2!c��눊S�Sj/Bb4ھ�SE�:�;�,�ar�j����3��eJ��$��B��
PR��6��x�S�c�$�_�u�Qd��@Z]W�B��B��~�+/S������e���5D�^\��H����<<����0uL�S��S����N=�8j��[Qߑ�a���s2��
E��O�FS�9<s��+`�m���;�4�]��f�
G6��J�U�QՔ�I�3$�ϓ*|sMŇ�� ��9�{���y�L�hGRC��l��+��%��/�Z��)/T|�:P��2�j������B�@Rأ�SZ�ԕ?S����?��x0u�(�iKGt�K�DVgi�b�����MIŉ�wA��z1Q�c��N;�E��T[�h�cR�i}:l�c���.�PF��v����ĊJ�����i���M��1u�管GPٕ�d#F�,Ԍ�������Qrޕ҄ �x�ԧW��0��s���,[c�.\.*��f
��7�K�����9�l�@���jzQɨѲ) v����1U���l@�����.��ӱ�!���bkWH�ש����@bC���\�_~0u�j��0N=�c���b�m˳�����"=H��1P�Uw����S�`���=��_}F�wsr�O:���LQ�ԩ�T�C��ɾ��\u�"`�%Z0���E�k���>�}�)���$I�9�p
�)���G�0��>�0u�����卜,�+�+u��»(��1u�*�n��V*��jy���s������q����D+�K3��RO��i�
��
�.����d��i>\���ԥ0���{@q�a�m\�ӽ��T����T����ԥ0u�iy�
K�� �z6�f�bK�{�8y�ʕY����[��ີ�o*���!��OE�;�F�9���t��u�i��9���O�������7Ri@�X�P���@ۙ��Y��I?��]��D�?�6��B���gC�Ji-���󯸒��͛����$���n��AD֭��L^!wډ�H��V
ƣ���1�+��1u�x�z���9���ΞI._��E���*^�P��e_�a�D���ެ��r�X�G�o��*sF�� &2��M��z$�ZÂ�S�B?v)�O��^�k���y#�|g���ґxͦ4+������N�s�[(e@�\��N%ωgH���H�Mķ���/W��:�Wv���~�n�����L�h��vjy��4#��R��cHk��)�f�
�����ұ�A 4���|6�;�Z�[�~������c���鏑��!dJv��S�a�&I_B�V>Z��Ag혷�Hz��\��gҝ2�l�l��rY��6�DqL=q�Z������'$��d��S�/Q~�Di��־�`q�j/<MR����:�v�v�� ��d�[����-���K[q����0�?&+��(�^4u�nL�S�uc�Fݘz�Q7�^�ԍ�'uc�Hݘz�R����T��z�.��;u=L����1�Vu�I{�;�*6Lp,jԁ��)����j<V�m5��۸�����#mI�����B���¾�e�]/ U���P�u�)��=j���TT����#=KJ�D:��k8ESe�f*lL��.���\"�z�W��ii����[!�*��>K�Q�\G�@��?��w_Q���{��*��խ%۶;J׃�17�}�=Unm� ��Zw�p*�z��l��a�x�52��T�u�3��u�]K(>��L^)[�o�]L$�Л����{��|�*9�2Ip@U�:<��8&��^:V�I�BǮ�Tl�z��a�| �:�n����M0ud�|�w�N�=�$��Z��!�ŋ��=���?�*�F�N*fL}k
��6%�b�����7uc�Fݘz�nd
��{b�6K��v�bD�v���4�ݸqэ��8cQѡG���&���K�в�?f̔(��[�vT�!1f�y�dE��Q���{��2#��i璽G/�3��z���.ٶ��h���h��#)S��K�E����]��{�C¶���0����0�)_��SU)~�	bE6y�E�z��� ���Evİ�p&A}����x���R��Ա2��Mz�`D6�m
*����-��ي����5{�Ǎ4����*����=�^---���u�u{��G,62c7Mf��5k��/�f6�l�Ъ�V�6�`��ז'�>��-A�u|�ot��������"���Zfb+f�R�y�S}���jc���ל9 � &�عQ��E��w���i�9�$��-�e[,�.�[��o)���5L�^��>3�t}�Ls��
J���EQ�.I�V�䲍v,����m�w֏�bҮ�1c[D��.��{'�+�&ב#��sY��*�:u�C*�u̹�����^bB�،18��G�.���1�R��)�N��
�N3��R2N`�:�L-�=);�{��7��z�*qѝBki&��w'3��m�(�����(�lޟL��qX�$�=xC��|Av�T�P�c����S⇳�l]L�ҳe�0u^ �P��px�K���S�_�L΃����C����Xt�NpcR��ߟ)�:u�cj��G�'��3U�%[9�]VL�Q�ש7����{�zfa{m��MEE]S��un�L�
�M�tL�ː����z!�oS/V*~L��L`T�����+rD����	ff�>_��6�V��jS�7�!0u$i۽9�S�h$U�]�9�Ի�s�SL��P��>߽߻�#Ҥt����~��g�BB���L���χO��:?�d�	�^E�?.�S�;�OR�؋(ƌ1k9�ԋ��1��|,�I�8A>��c{��n����E�ϒ�ܶ�w��q�Sٵ�u�pjy���b�9!�luY	�)?��|L��K�P���|��ǹ��o�|=�tꮲEF3E�I�!G��u�1dvy�&�cL��{���[���	2�3/"�r>��_�_��'�[}�����o���ӏ�|L%%�2'i�Q"=[B�.R�5\n��~#��ڸ�z�T���oPəP�yW
Ό���>_��ߧl���c����a*#R?�3F'0Yr/�Q�������N�N�*)����s��gDH�˃-�?@~�\�K���RP���`�9��\�ceVچ�ъ��Jm0f�~�Y��J��~?�H����Df�z<'�(�n���.�r��v�y[���u��_���#�K���'���R��wKv_���H*f�(��|5�L���L8G1E�e���|(�uS/�S7L,�.K�S�"�V=8���͑��0>�k�C�)0�m�ﲛ���A[
�0�c�����0#N�"�kbǰ�_`S`�R\���2�B�0��"���\���3��ٗ��u̐��:Ì�k$1�-��)0uC��2^��3!�f5L�F�^�}����m.3"���5�_�� C�m*L�C�X)��G
�{�<���ѩ�o��0��&���3�K�OVP���*����1��6U��t�e�9�oc��͂���3{�'����/6z������=����Aw����/���o Y6��װ#���u��G�z�i�kxg�_�}��y�<bS�4r�;R)I�,����W�z�뗗�C��QiwW�`�_�����?YH�N?Z�n�5��gk3�[�G埚�{�-�u�a��,��U8@��3��R���>`�jh��o��5�uH?��������.[������}�}�����y��oPൗ%�C.��/�R��-����ﭯ���E<Ss�T����ڥ�;��*L!t����m�G� �2��hż��� �s�G�|�~�'q����io"��F�e?H�0�'��z�9䠴�cu`�L�a��|̡���|\t�b�(Oc�}3%Ķl;��B�j���0^����r�J�C��a_��~�ɴ�1uMDW٘�*�!�/)�q
՞u���޾��/pi�4me���y�5=)�v��F�{I�M����� � �i�m���M~g��y�*� �_Pt�JR ���@:җ�U���ܐ��(��	U�ȿ)���4u����;tk���3Y<K� ��N�V�~�߱M7�A`F�'������e�ЕǘA8 H�4�(�aJ
3FS&��8a�].	�:�8�o�J��H���_������P��L]
9��<Q[x��GW,��w_']���_}.T�?R݅���#a�01�����l����kfH���콕����N%װ�0�J
<�$y7�eSw�Sl�m��ʙ����㟤uF��Ϥ���	�"^C��撰_����� ���.n�1)� �/R6����P���ҭۇM�{H�lslbL=�� D���_��z~Y��V�Kv�&�^Aq�ϴ~��%9�P������uR~�A=T!4��=�-�(�z�fݠ�W%~�q�A>��c�I#���i@�*(�5���H�x����S���H~��sB�_򞸍�=X3�M�C8��8�r�(ژu�EH�h���T҂���\���PAb�e*XL��L���w�1�?��MS�1�nʖ�����<�c�s�[    IEND�B`�PK   �p1Y�?HU!  B#  /   images/585092fd-6de4-462f-8499-92296fb2c536.png�U�S��]:��n���	i�F�;�F:�����n���n�x����	�;s�ܹ����=s�<��@lJl   TT���� $lL��m�����EA� ���o#��hB�]R���u�~�t�0q� xxx��8ڹ��|����l�y*A	 0�+ʂ5=�N�<5g��=k�K��"3c�����s�zhj>����v8�*����U�]635����D2a���Dc������M�P~��"z3����l�Μ�ws�+<����1v��2nh���0�*�� �dz�̗.�`;7)�G�fK{�"j�R��6G��e��o���<��Z��o5І�h��+u�8oi~�'�f;- C9p�]t���F�,��0^M1��D�K��7T��*��F&���Jb��{.����a���"�P�R�9)��H��G��3qx�N��
����=��Sp�IP���=YQ#��Q-��\F�A� /R}cЩs�@} 1���H%��4�k��(6K
w�Uxt��c��[?2
��Gh 6P_�-���(�QXA1��+6o����ws��p�&E�{�Y�X��"�UPӊr�K��=1��8��K�K o��H�hV����[9�p~S��}wuZC�p=3��GPZ�d��-��jn7��~�ʸ���O�֜�����3iZ]2nT�p�'/��g�}�iU*�k�u��V��gOaG���:p�r�N�@��^\��	^������N��ś���4��Q���S��g�S4O_��&�\k����ീ�A촱4��N��u3k&lE�&K��q!� C؁HsCY��ۆ�@�[<�I����|�h5�@w��6�:<��#�w�\�ն�iI�m��G������,�}�f�ԁq�cc}�zu���'�4�6@[�KW���<��T����4.IōˍY�*��1�ف�+���R	^��>�]Ư�;W��d���tV5��C�xłyx�^hE�윽���d���7��7�S�+tP2�]��1��E�9��j����60��Aʗ}�e��3�vi#�k�cNv���� M�U����D�@E���y�̴o�U�;�]�t��n(-�"�B�}�2v?e���}�;�{��'��{�A�/7J�3�f�#��{2���t7�0����-��'@~z������
 K[���ϗYSIܯ�K�>���@ �p�^��z�k�w}�}���f�,��sT�yzU͑6�3s�7G@k��1u���ˀ�k7��q�������������>տ^���� ݔƥC��,U:V��3]�u�������&C��j!���W�>ȹ���/be\~Ii
�l+�����`$E����Χ�"����O*������|䢤W����'mo����
��glFE��_$�)�xK�EC�~H"/לiVcƁ.��4��tFNX�/��Z�3���Tlڶ��đ�Q�"F�VV��ե<_Z��������X�>��ADr�_��-��2�M��[���Y�£����R�"����R����}�$�b�E��x�@#���H>g� B�ӆ�z��F�\��@tR�>��d���9�����8������N�1~��Յ�ly�H*�n(�d5��cؑLG�s3����j=m��� 0��R�ˋT�eM�-֨�B.u&o]��?,��aGYA��i�L�s�x!�5�7�������hpy*-�l�_�FӹaQB��s��c��ٍ��4?��\�uO��`�j�!�����|*����P�嵙�1�@m�º�t�:���g(�<g�3�=��u&?�[GG �ڗ���#�ڐ4�Я)ٯ.���wޅ����0����(-�A����yC�>[}5||���[�
}	~�6T�J���9��x�x�4DE�|��_.�1�.��l�6�Gtj��;o}B��@�����̛��/R��J�q
!3�j0���[@2���}8Cv��\�MV�iM�(�L���� �G/�~S�߳����������~"���
������ߋ5�yW�O�c�2|*��[���3j.-��ބ�"���rmʅ��m����߈dd��$NQP���f�546	{���|wRZ�I)/��Pάk$�3�6����~�RfU������u�ס��R��tT�6�u��S#����zd��y�w^�Y��E�'�����H`��i�1�"+�ˍW����	��W��0r䳒s~�tC��5�n�kZ:f-��j�7��g�q����7��#M|�<����
�梕ѭ����+�E}#
�̸sૃQ�z�� Q[o�伿��:!�ޗ�qꏳL���XY��p;~��~���ΩEMBD�sw�M�!-�j8�Y��dT��k���4	����c�*[��P�4�4�.����
�o���� ����x��t��������ye�o+w��T�g��}c�;�#<�H�<geζ�����_S��R��5pVSP��{���p��7�n��P��<)�ͷH:��uj�RAҦ�(�����ݳ��/eB=�g=v�	�U���62#]75Gd��nt|l��s+��hfn�ɥ�M�N�Om�"�aTF�'?֖旱.��|H"�ǚ����ϛ�>lس�r��L���޷7	!�`US=�>4�煖W�FNú��(q�asǟ�Tc��6P����Ie���1�S"��T.���n7u!�f4����os{kW����/w*�����.��%&�b>�p%�ݾ�%ߌ���W�'����q���O�Qf�B��!n8�sn
�~j~���|7�VU�Wj;CH��99��v��\QA���o�;�S�lj�٪V��Wf4��H2�8��د38�T����ėh#�f[����M@�E�'4�Yu޹�������e��7�e�ٞ�2v�+���?=��9)��Q�#�S=Bxo�k�0֔��2��l�M'}��B�r_�f��{�7~�W����<|KD��-C�4��Uʼ�jHa�
m����ث8��N\����ZS���Vڋ��G���瞾��l��zn����'��l;�W�m�K8G	���[��?�c>H���J0�c�����;�?��w�6g��2��(�1AQ���M�y���[�d��T@�i�-����X[X�B���f�0G�k�d�_��7w���1F<�l]�>�^��M�	��q����H�KzmY�82�#�s廛��E>.&�۳�ǥ�g0c&,h���6u*����U!��2J�|^Q����9:gr�x����]-�*o�F�̱�`��E�@�Jho1N�2[�^S���Zf�:?�t���T�Řl!\X�����
�0hP�"�w{ɭ��RiDc ;a8Ir���f�[��}�o"P�'��OG&$~��4��|nj�2��oǺ��Ye��!�<?��KY�:5�+f
���ɡ�8��\����L�����/
G�C��Բ�9%vJ������X������E���7VR/A*��sBN`L�p9#�(�9���c�J 9�O����FOY��a��k�IƘ�����BpBSLI�*׷�G&��gL�a��J� .�rǥ�6�.v�_mO{拃��~_�,�a��y6��@��4m�\6���B_�	L�𣖏���g�֜疸�TüO}�>�㇁���������>��	o<ƍ�������>�x3���H��Z;�)x��t���v��h䏲�Ws��ѣM�JgBSW׻/{=�6Y�/}�G�a�|Tၸ[3��9ހD�)l��?M�7�\ա��6���]fq�;�|�0@	�/L�IZS^|�a%��Vz�����9i���G���﷞�;5o��.p����7�X`GD`t>�-�Y���0��o���h�p3��r��;z�q�����B���^�����`�vH�%�%ͭv(x��X}�c;����}`����H��yL>0�`��m���[0g��W�� )Fr�Sf�$m[Kx��z�	�۫�G%�R�O��
J��+��F�]v4�9���;I����L���8��ҍ���wN)i1j���c�T&�M"l�"��L7�7���)=\� ����z�g�a��L*t�jB�g'�:2���������2Оt�raȧR��y����8��YP�Oh���a$6�!8n����,?��C'���.�M��#����nj� �~��K�nA�;�k�u�/@G�]S(�<k�lZ��Go��Ϊ��\c�e%�d��k�1i�"�5� ��=��t?���@��ƕ�8v���wE�Y������h*����r:Ɯ?�ms����l�Rx���~���o����~�F	�cں�?�Q�U
!t�����mEE�5qs��u���2�Y���-IJ���<��&�KC�B2���ʀ�]~*IQ�%.�Q>9w+3�@^�L]���`@X4���r�Æ{2�`)��<>nLʾ�Bk0<;���yK����ޘ�J5�A����n������HƗkh�K	�%,�û��Y�K�>�b����T�֓�P� � �ΨR�V���fM�{��;/q,T ���5m��'3��6s�׼o���a�֯b-x�#��}�q�Kv�7i�O��R?@Ӣp���/'e޺"�X��ɏ�����	-�*�p%����A���
�����?��nD��@�\�f�t���7n������XϘ��h_I�ˣ�1!^hf|�VS����.�'+�?߀>��^AP�fg��w��1!蘧qs�����xAp?�Ы�㽋��`z����6�'���f:�8��l@�
˺R��l�@<*���h7�Z���<Xy�{�#���L%�v'S~W��z��T9O���gc���k�U3�@�#���U�z����WAV����S��om�:Gx����U���xEf��b�J��:��,�D���������_��a��N�(����ο^^2l����j]�������#��Z,��^t�x��&x����%�A�9W�"�{~v}����t.�����H��$�h[o_#�fá�<�,��X?hr�x�IȮPJ�n�w�����d�&�(x��L�����K��^�BQ��lc-$����mog��v��>F���}�|�S}g(n�y,�\e��C}uv�i.u�����~Rm�*��MÀ[�9Va�/��T�ę�M��0�fz�ȁ�����E<��??��3�N�+fk%�5z
?�#f�(�*�����z��'�EH�
�:pơ���3tL-�?� ףg�Y	�h�wq3�wY��Ë�R\�d�{�����c{|���㄂<����/S��Y���f������,��C_�Y���Sm���ay��.cy`�n�͘����!Z*L݌����63�us3ˣ�c ��ݵ�h�~C%�A-�.�&��`Ƀi�U�H�*�~r,��i�'a����ӂ�����k,eFJ�`w�5o+���D|d�ɰ�KP��d�:M�`q��~���H�@K�y��@� �cidf�_�=c��`�b�yJ��-O�8k}��b}x@���Qr�bIi�\P3��,�a�!�_s�����K<����v�y;��j�WU�4 {��}N�b��&�$dL8�[c
������*�ܙ�8�B#F4�F$��*�~ᚾ>�IL��D\��7�6y�lHY�E��C)3%�᝶�nzl��ë&�G�$&Փ�B���'�`l *#��͙G��i�7dij�ߟ36�Fs��e
��xW�<Jj�i�y��꣰`\�H��b$����;�c�V��DRŷ	��\U��ͭ��y�آÚ,x�{��K��R?��E %�GU���:i�@Z�H�������٥�o�r������p��9m84!��9��q�P;���c������q�N���`�<�_m�_-�O�}�w\�N�Z6���ƾ�M��՞�������Dٙ�b/�BW�M�XT�8�y�����8CKі���8�h���T/\T
O�Z�V�L=��x���,��x�v����J%D�����i��[]^,��G�����>z�I1�E����'[�4kq����((fܒk�x�`�9�Ń�7⏑�Z/t1�$W���{�t��s���ܠ�UO�s"i���'�X3���>2�������O��j�#�]!���IhJ�D<]���������I�81��2��6�|q�iǂ<���Nr��;9w�=������8,�X�&p`	��9w\
VG.�8.q�EM�iY���@��q�1m�j߅6�}�	��Q��su��`�w�Q�i�[�l�!fg�>��m���wM$D^��+|>:��˖ޫ��Yߝ.6K�=0č�ө��e���h�s�{���x\��Y���*�f����\r.�
DQy:���[t(5�jM���d$���K� l#5�wǐ!��ɿ��Y��D*��;!��!9�wŲ)��
]�Q	�ֿ�/��q���������!H6���U�o>1��A*CP|�g����)v�J�������~A.-�rE�6.�(����$.���H�)�#t�U��+� �G����_��?���/�~��fO��)|rn~���S�Fo�7���R5��|���:�?N�d��b���g*-J�[�'ʺΝ�V���0��KӠ��K&H�'�������V����!��rC����ڳ˸��|5i�r$KȳA$��r�h�P�-T�'z�g��@�H`�;�<)�E�>��%^�H�6����n�����M���r�\�h}�*��V�4��Q�	����G������AR�M��G!N����v/0�����zy�����Q�!�WNqY
��o�04m�[�9�qQp��o�W�fSB(Ku��#�<'��'ϭ��gB�_0pA�bٝݪW�FX�l��I��N���2�&�?�����0(�P����=]D[�>302lv��̫��<⍌�^¤��q�Z�О���Jі�H�⿷~��[>�U�R lļ�R$y��!*�(ǻa@}Ne��`&<�!�I�ʐ���ć��m����+�&@�E'Hz9b�o&�R���&-�v�hyA��<�}B���Ҥg�(�!�%�jCP!G�jNnnD���ژd���.Π�i�U7L����\[���	.����!�A�{ Q�Y��?m��ak��f�1.00�S��!�sSA��f�%�Np��(�����-<��t�d ��0���	j�$L;j��
�\�p���ڱ�������{#8�x�ˌjN�TnU��f4��u�o�9�uD����F<R��e~�>�Kb���$3���D��x�漹��h��x4��a@������_Fc-�(��7���O h?��~I+6�~��/���h�Y�i��_�A	�������eT�$Ўl�U�3:
U:�P��W�6=��8K�V��7yѰ�*��$C�O�d�J�D-��M�S>EKN�*%Y9*�B絥���*7'n�JI`�CFʄ�w�����	C�:�.WP��1%�3	�[�lC�V��G�;�h�Pd��]4G���P��l4�=@��2����?�#N��µ��F��!_�Sm�4����dY���+w��V�r;�Ovd=X�~ɠd�3(,�WtL�jG|��/�B>�Gi}%聖3�1�T`~�#$���I��a��AN�'���,|bHM�3�-�"_�_4��1|���P��8E����,�@J��X*[)<߁�2���r��B�¼#�a�=�%ە��A�Wߝݷ8�^F7�fz��R�b�M�n-�k�A��\t��_P՜~f�MG'�sg������Rn�7�Ѻ����"��6�5�;(���~A�nԹ�
���s��6ݑ�����Z&� ���c�I�y�?�l����ђA$�͟��9ȧ���f��cPUg��	(u�>#
㏾��	gA̡ɁX΄ZcX.砮���hT~Q�v�z#���ph��'7��Z��Y��Z"��Y���b��p��2�s����hS5/W���G�h
=�=ZY5'���4��3�����WY'�����,Cf����d�:���*���#�W%��W�x�s��_U�I�홗�����1\)�e�Er,s5�r��YH�H�q�1û��@2D�R6���
�6y`jWDA2+9���Kf�L��9l.LU��v.�@�����x����X��񪼗c��`2�(	�N/΁����΃B�,��F9S8m[����Jq[�07w,+��
zE>�M@}����V� K�ZspK�	�щ����M݈�D�-MiuQ�|g�9{ٝ��|�C�o�k�n��Xdy*@��*m�����R�g�1R-Ks���9�d��j=s1�m��x�sms�O�1��[��Te+!�A�PK   �p1Y(-�� 3S /   images/a48cfa0d-8c50-4ef1-a8da-0cf94db079c2.png�{�?��wT�]��V�U��Mk�A��wmj���FԮZ�j׊[����=k$���\z�����_��W".����>�u��TW���K����k�@W&@ ���ȀO��D�˞O�t����~�|�M��bn��&iv��>���{��j������p>'O+K7>W���]�H��]���Iߏ&z��ޜ����uJ�{O_<}z�^��;2&]�IZ&��-�>�{=?��@>���|�;�Q�}9E�3�7��Bu?��c}�����J�G��~�i�4�_�����V�&<Uwb����l�]���w*I�}?s������!����Y��w}������寂��]"��R�Ƴ+�wy�ܞ��{>�K&r�'��x���(��`��� Ktg��Rc�{�����؛��8�fV��;�Sy2��ͅ�H��
wp~Ȩmns�1hl��8�����#�����.��x?�d��'��������Y�������@vA��{�[D�	i���.��]�W�bU�GĐ�N!�Ch/��i�"��M��n�P^�$�󆶒B����C��sM����|>�!^����Qbȴ]v&@�w/�
��ܚ�8����?!�J�=x�@W�L�?S/���j���AN	Z]��˨zւ���f���C��>K�p�c�V^��%����"���X��8.���p�j�䟋�~ZX��w��uF�%��Qrz	_���{ ,e�פ?���c��#��`�j�	�Ŧ��`�ӯ�C.ӏ� ��W��yr���Q��N�9w)à�>O�Tu*�Ƈ��G{���3��z	#M��ɷb�^��Q����ٺ�}	_��$|n��fU����ǐ|X����{|j��x_A2b�P1_�ղ,��y6ʏ$��е s�-��8���&YQM��?k7z�u�� ;C��2W�с��^=�ᇂ+���2�C��W+#ْ�%��,p$�3�iv��9�^S�3��쪹B�G���t���:%F��N�e��+�T�4���c�3��iD�����ٸ�$��+amEM����z���� �b���aq�䢸ކ�@S�y�������-i`�d�h� z�����}t5b]�#�)�gݼĳr0��x�\-G߿Ly��0x����̋	�����������Ff�L���d|��k��
���/_���[�����M䪙�PMY�(oM���h~ڔ��X3��,mc�M�� �Z%�k��p�K����w����M�N:���'	wt��eVQf�g�|�߷��|Z䘢]���d9I�i�#sa�o����S�QF-�ٛ�n�Qp<��9��F�n�����OX,���Y���({������h�[Ɍ���!�}+pK܋�o���t��h��(J�1�9��i��jcu�i�l2�ϫB���+d�e[o2E5M,�W^�s�>��K�
��3jX���si������[BP��n���>a�\���pN���Z�CP���.�q�[|�3(,��6�e݊U.g�M� �S�.�_q3O��<���U�Y�Ǹ�D���@�hg~@�H�o7X�o{�.���A[5�민0���)˿�/�>��f� Zc�OBW��������o����;��ug�ܽC^��UkF 9!����Ɲ:7h������\�}�kF�_�I ����� C0��¿E(d%xA���$ZG�C����m[�j��`N|qӿ��,0K�֣�x�Ⱦo6}ȷ���Y������8Cb����ʚ���m��ǉ|i��-����
�����(Uش?u��O l��_-?-��GY�I;c�x`m^8z����������JV644쑼��h�S8>����#���e��U�&I�&�x_=���?С�\����7Z�_�����Q����a1>��q�꿸[S���''E���''������[����?QP�;�̇�}R�
��8<�Z'��`ó�r�T�f�/%����K��m�/y���3�N�u���?�;��m�g�,������=8�N�ѐʐ9��+>��ose������đxF'@=}���]��C�������4x��i���y��6k!ᮓ�}Q�:��-�s�?�̵�P2/j*[������_�����p��g]Ɯ�ZX��T�]w¥8��#����D��t�
�Ӛ��(Q���l��сh������=���ɹj���x�(#���MM��}�U�^Vq,��j"Dd��G�7D������ �a�`!�*
~㯛%z�Y֮�i�s{$5I���$蠅VH�i�s!�J�U�~O�[y?�ͯԒ��8�H�B�Z�=ԥ�$�z4�/ơ= t-_;=C=�S�+)���z�}�O�}���|�O����l�.e4��u����d��,�.Ã���i��\�u�����!A�d)�g@d��.��x�$��T���O�x��n�����o������F�y�^f��ip�Ñ � {�/��n��m�����c�ծ��uߎsL���&V)b�B�#�(s~;h�h�/W��z��S5�5����+WO�"��l>K��ux��5�W*�;G$���S��iv��5w�?R�w<����� |⺑�B�G(�T)�!�;|cn0�<Hמ�����ɂF]��Z���-!	Tx�������2�Ds�l���w����J=	������?��6�T�ڃ���xG)�P������G�����: -���!Hw�Zho�I9�^#�����8�4Z3�r6��/�z�s�i��"<۟s��}J�|�rk������|�C<Bkj˩H�3�+��:[2�/�I��[���}��4��Ӿ����9���i���T8�>{Q��R��/-�]�
����G�<����q���q�(ry�fY^����7�uroԵ�-�8~���P���}��h2�[<�9����̞�z>.4����[��?�bf�
�-��SK������QN�W'�↪.i�ǯ���-�� ԓ[�����ݺf�^�\��������m2��a������aj���cs�Ԡ���;
ې�YQ��ۋ��O��ޕ� s%K�����=�J�f|�v������_�V�'���Gq܆�Z_��� yޥ?�7~q��T�VSsf��p��l#w����w����]�c1)�n�s6��S	OW�F�0���߅\�2��Gu�g~����x��Ʃ+]%#4m�����<Ϫ�a�O��LΘO�Žp�ҳ�R�#�n32�8�"��8��t����^�)u��DS�\��`>Lǝf�����+1;4�.�~	fg<��tɋA4_��^�zU�ؘ���$�zJ�=8	��/��j7Е*�u���0��������Z<>mV����:b�Qk�]L��G��#��+�<� �m�+���s^q�6�}����&����;�	u3�d�"��˙��z裠�+����szZ����r��#����&jm�sOf�Gܢ7�GĿ��z^<��k�۝���zW�d���l��l��th�z�TƷb9�O0�D�y���tF�B�#]�p�y�
BVx���Ŋ*L1���$�4�[W�a���8��g˯ښb`��ܔs�Y��9�Eڷx�m $!Hů<F��ٕ��'!b�#�:�ޠ����ז�d;�y�N�Z�E-�1�ğ2;��1{��^���7	v�A�w�xj���L=1���㺝�R�Q��\O�4�b�C�]K0��/�����2IE��(L���֫���j��#�n��6rh�������@7��ə�n�z�V�qŀ��O\����,�r�}o��\w`�%�E��\�
��σ��jcz��.`�ބ_�Ǵ?�B��-��>�0���fI ��۩j8��Ýc�4����;��нtT�JKN��#��Y����vc��&&C���,:}2'�Y^�¾D�@�_N�ù�+PF�6�na�!�O�y������%^�Z��(�1�hk���(p�d��5�����2��p�>(	�m+��uL Y�[�&���& �F��evx�Ķ�q���uL���W�oo�Ȃ�����3y�I��=�Ho>���l������]�n�NK��0]W�*B�|����pA�w��s���<_�|GA�{1��&:�O;��֟(�o��L�,�����W'W���+����\)[0���|.A��k�����\���sx޶�_�B\��+N@M�i����w�W�XeO�8[���fD.��N�$�oͥ���Vo�{!�����tsN��nJ۾���"E�ʥ�+1�KG�Q��?g�д0-��>��[G�W��<}�6jQ���w�P��:W��	��	c=���z��%Ƅ�߷���h���jt�K9ǝI�u��5�q'f��Z�I�ta�f/�<V�$����۷��8��XYW�~�3�>�R*3X��������]7v)c��`J��j^g��D'�^[�A��T�m7|!^�')^��7>Ԗ�{����:	�����q�DU�&���-Ju�_ByKc�%�~ٶ�McF����'�3���%_�(#6=��%�\��@_Л8!�;;N�[�q8Pp� �CtS,L	;�U|��)/�=^$v~��N҇%`c�*�{[���xS�覠|id�Cl�C�R6�9��<I@�Y�s��(#g���^��:j�W�̯㴮���N�cO��<;� ��&����0�Z���20;���Wt[~m\п1y�����)�C�+���S�g:A�A�~�0Vg�~�`�q��n��'�N�P���k���V�~6��D���T�� ���gQ�$��2}1�ǒ��O��թ%��%_�F,_3,�ֺ�ά8��ٓ*������k�N�z��"��k�~l9��u�E51�p�X�\D��SUl�K��zy��Q���hb%���&&�� �h�-��5���i�u�+Ħ���boiD�Eޢ'^�/0�e6/�����	����0㢅9��윔��^U�	C��k��5�{'d
`�t�q��/=��N������\��۞���v��G��X�����	TS��?�ܭd�$v)IK�O�Ň��9�;&>\�	�1,�U�.c�.{�LT�-_�5����V�m��
�1��{�kr�ls��P<9'*�do=?.Jy�d���pt �!��Z�]9��lƿ�����ټ5s�q�mT�$�0E?yo��Y����kcRY�7��t9W�������&��+��ʞk�Ki� �4:�?z���)+�#��	{m5�������]i�l8k�/�-WҦ;��|p F��z�4��`r/�`���j���T�(���F#�`�]Z����J�X�[#�t&V�j�9���}��go���s~�b<���nqc���jVb8p��*��/�(�"{Ӊ�.�i���sQ��5!�qܴ�Li�^-E]��1�D��ȣ���|�W��c��4m[���ObB�aJ�~{aFȏ0��lᨾ�JylW�cfГ��|������.\R1��2��'B�����|7c��ǋ�z��N�PU���K7�}�����V
Z�-�yG�������{�������T̛���!+�_ǜ�&�Ҭ��B�����E������>�z9ꃇNEK�g?���5�@���v�Fh�s���)�X;�W>>l���<�w�l�Mjx}��Tv�w�WkAħp5��J�=�ԕ^l5�$�
̮����#m'����{T�{�{I7s�~�䕁QH��9�)�%�1�g�4��
<��.J	u%�o�qջ6�:���e/ �)�K�M*��b�uE]�hD��g�K�Xt���`��[�a������V=F�[���l�V��0O����fT��*�=U^���!9n����{0C�.?X�'ivK8a��gi��z����.T>�d$�*Ε8�za%32V�����Fze���������c?ߞT7��Qn���Y�lt�.�@3(��:Z��2�����LI(��#�
�q���u�e,rk)��-��hK�l��)�G~� Q������;�H=qH����yǺP--��no���>�'��F�P��
}g�#�L�tZ���h�J�o0]>�h�r���׳�4{0�M.�q�̲¿��|3��@���8A1�q�}ذ.���|sͼ�S\�f	?WU��3�a��6_I+����ƣ����Y�n)U�=LCkJ���~�]�(u=�p�b�������W9k�Ntʮ�,�2(�G�m0�Ă�S�흥;a�S�5Uk���X�L_�4�A��x��ђXk� ���4�.��n���G�_̭�=m��Ov[\�%:�?<~@]|�ʹ�s/2��(�Nɗ���*m@� �[��>4���� ˿�-(4�!w)
#'��S%'hλ�������Vr>�� �������w�v�!��!U����de�NW�7��zP��-�U�B��{�_��F��p�?l�˜شo�.�FA�82�ةq�K �7�E����nz�S����5'���O�as���;+��SG���E(�+�i[��_�I��v�S��Ş	�Nh)h�S+e+��C$ȴ���v�fmHo#*-t$�ِͨ`��M�x���[��P�\h�>u�d�ߤ*���9���@e}�����5!V�[֟���C5&�ʗO��Y�J|���M ��̺�Kىy� ��z�0�s�׽Zyx�A&>M�jS�1f�p6�3dKW��a?��U/]S:(���͛��_�G�l�*������4(\�9_h�U���@��QS���M�&���;��??����Ź�+�	Y��ܤn�a��_5���\�W
��)���V�_����F�EK�v2�����͉U8t��ݗ�W��$��,T�T����x@��t��?<�^}�S��}Mx�_��B�h�&_�PŢ��G�Е��glV7S+4�����6+�C��CJ�3,n���y&g�q��+�6�b���eQeq"*K"8S�U��U^^4j�:<�����I�_[O׫�V�b���	th�Ac����7�l��T6��B��,���,����L�=�:�=�fO?�7j^��*��ν����)D3������(~��Da����b��5�v� XY�	�7��qR��Jv�bP1��<����FDV���Q�_���԰`è6�;���B�j�j����M�Op�+�&ۆ�(�:<����6w}9���wЬ��~�hiX�Q���G<3Hvi{&�2Y{�y�^w^2�ސ�C-÷J`�19�V��ީ$u�{�J����D�kQ��# d���VSAtA�c�K���P���XdR�V��=H�2Y�*�]�>���f�����4:'{Dlt(�����B�+hO��}5ƀ��z�MkqZ��߼�`R��lQ�G�̽(��0�P�DZ�mt�����]�}韓l�����9+*� iX@�XY@'`�y~*P���d��ޢW�C����a`ҩ�;:��9Y����A�^�o�����ɻ�����Y̛�yî�d�/S���,.����O��^��\��j#�+�z�� `���/X�,q�<�+�u�I��QBC�!�X��'	'�(�>���?���D�$�y���o�x옝;���R�����|9Bڙ����.g~r�B��ɺ+�u�N�]a�Ĭ=�[���Y��2��'�zQV�:憶�5�wi!��.�ܿ����*l�jS�u�1������Ϳ7D�Ž��Luw��H�OD�.n���A3�Λ�� Om.P'L=����@R�|6֧��y+��d��":��)%pd��И<�c`fVN��p���r�:��h��vsR�mY�g,�����-���⊮D��xR]�O�v=�c��8AY��NeҰo�*�5�r��#�~�_��[��=�p�_��[S� ��/Tr�T�40���M�؛�_�
dOv��tzEykL=8�Ňe�ؾ��:U\%�[��rs�'� �?=
cE^�,�-�+�W_��\���d��3�B�*G�T�'OH%s׊�ǵ��͞)0;�I��IrAB�Bu����N��L�y$s��S�{j������#n!��6{,���F�D��c�}�Ԙ�-���IZ�K�]�0�,��lz۾}�xF�l��Z\�N��jB�2�^�P_�)�8�DH��t`���h{kv�{'�d��~*���ٮ��w���w3�CJx��qDv����WPB�E�`�9��.stѬ`9��D��Boު�-;�o�2�Xȿ_RCz��?4��V�2<����U"&t�QH����(���YC*9�x�J�lx�p�#��Hj�%=}�U�*W~S���i�M�v���Z1�M*I1r�	��Ȳ�_,�+.�/��hf����;Fc{�����G	$ U�}gNV���b H���y�W��@�vF�,���@��e�͡,y p���d�L� �i���C�hd��|[n�!�i�Q��
�(xp��{���q&`}�wĠy��l�4�jB�>�M�3��2T��E@�a�=�طѦ9��y�v�6��X�b�~qI5S-�
ğB\/L�\�l�3ڇ��\�~��g��ߜW����FJ̧�u�]œ��}5�u�?�c�#������!�	L"{K�?.�>���k��%�8�g��Wn�,Y����3g%G��g`V�����}���S�A9kx���c?�M�e_X���0;����|"���~�j�łƸ�*Xo�Jiɧ'��9;S�'�r���ާ�F��*%4�i|��D��'�CCb FV�7��S�s)8��k����X�~'!�XX[�"q�PtBK�8t��u������{y�bԌτ�9nK�oړj����S����� w�B)��R|��}�L|[�(�5�K_�1�N�)c��v5����ڥd��M���z��wa����ə�bD\Dx���Ѕ��8 ������[�0����]�}�����˩�����K��?؋����66�쯩K-� 	��qW�9�G/<1�e׬����x�u
��5�;��;�nST��9�f��
� ��_������~Z7.��/��}�ԧ~;ҤM_��[������5Ɉ�cր�v��i�e��H���<V
UԬ�&�*����e�6uA|U2��Љ�2�ߠ�"����2F�d�g�*�RM@:b�vʽOV ���/�[W�G�$f-���V�Q�����l�ӷ{�����NA���X����4u� �����'3����ee��'�@���u	��$'F7��ڸ�4'v��K�Bm��A��1���.��i�c0%��RKN\6ȏ͏l)Y���D:Ӑ�<8�-�ey��]T�z}����[���Y�{���#g�J���e�~�&�������fL�1��P�`R����8(P������6��i ��N?-D���j8S�FtĽ�(�}�'˒�+����S�jUUUm{��v���¯l��6�h�;�☹�|�݋��G�Y�2�^�e�53H�6�ڔ�����)k�ɇ�y�lT[hUq"fb�)�)E���!'f.s�*�:��g�)�v ��ރ0���
��6�vY!0S�<�|�@(l��ɉu���˂#����>�"�.�&�T� �&�N���*ߋ�#Q�.�v����,n�ҋ�n�@DW��h��A�`?���r��8t�"�NE��(@�:uo�����Y�f	��n���qS;$¿�^���m����Es�"���h<k��)j�K�pfR��s��c.��J1~[5y�04����@ G�'��߷4K: '����[���<�n��j�/�ج������nz��(��GC������]c}��֜�@?��u+ؾ�X?�
h���Mk"�9�"��vG�4̹�� ��%�G���7�(���
��D
�,�&�d�/{"#DD
+�.5ԍ������e��>d��wc��Ƿ�D�E٥�m����|"f2عk��WJ�i���X��TG�?�`NZ%��Z�V*���]c��]���� P�_H?;,?��v��������4������vhT�k��``��F0IyN�ʩp1Z�V���q[?����p�e�BQQA�>J5��A����������d�������K� �H����AK����D�[ނ�H֡�:=��ќ�����r;!~�d�W�Jo,a3�6��e���ʏ��ؖ%  ����-M�O��V�{3�E��փ�&��5Y?�=��k|��"
�%ԥ�e��8�Q�do����6B�ݳ�s�{�nݹ:��1ݚ%�5��]��0�����9$Q� A�uy�Q}�%����L�~�v�*t��'mt���h��d�V��5�OF..鎻��T������d�6!Vw�mwݼM�s@��RZ����Qu�[�BSڏ�/VBn�%������k�L��yv�4�f�8y�>�dE�3���X��i)�듇��s����e��ү]�O�X���8��v'b���
��ս!��oLQ]���$@�;�0j�U{'�r�&�n�&��BB�m>�V�� �����n۵T8�w�Ԝ_#ߧ?Z���xT�
�$�]�f���k!��&�nY����צ�X� G�y��
�o��7��Nk=�S��g�6C'=����fAO).��/!y�n�\�x��|5s0O������ƺ_/_���-�`���4� z%�|_#P͓|�H��zDmu��W���rQ���X�k�Ut��,R���~���6w�B1"�醄��U����K>-p�RɽFA%2���n�5� ���5�v.s�? *tA�lˁ��v˗��2za�D.y��𨋛N��g�8P�E)맸i%�})��3�@Bz��sb����Ȣ2��L�M����#b@rZ�o�I�a��z � 	ur�i���˩}��2����,n,\�RA�ECGS���0�	QMM� �"��j*K�R��NE|Ŀ�?S,8)��~m	.yb�������~�A���fHוO�(A���:-,<7��"��'��x���4�t�u'�lȴ
��C+��mvȕ#<��Jv)��j{wm.B��	 �i��=D�00�W �k�Ut>7��i��)�o�d� �>��& {���KT��L����8鍇K�*;�8v �X��/9p
��]	�B5~�r�CJ�`�6"D�М��u�� �}L�DW0�0�t� ��4��|�&IP����hZPev;[��7�
�h�{�Yu|�`N�b~n@@��Ad�т���"�J'C^���\�]lI3j7�t[�ߩ$��Kٳ=�!�xM���va�4�6�ޟ��o���ϮS��B��]��4��qL������ȥ7��r�b�$ ��t�`�H�t���)A@�6���؝'J�@f��L��V�h#���nnG��|e�3hU�O{vY�]�E kI,�oM��lY݊4V0	G ��)���R"/��z��C���a`�b1b�/��iV�x�L�D�zF9����fu'���I��� 㿼j���Qs~6߻���"��k�=�nj�[��A�3T�I����=nzZv�VT$����>$G�(��8�A�t�N㲌���#�ep�����M;��j��5F��B$T��?	W���ڞG_�}+mˆ�~b.�Q�@ɟ���D��%hu��µG�z�q�Rڝ�����V�ZE�;�?��MU3P�JRz[��Rp�9�����w��I�?΅Tĵ�;F�A+��Y��,^��v�A1��uϵ�Q��>%)�����F.�Xo=%��>i
Ȳ0���fj>���\|��%�x�e�PG_��NWW*`��3��\꬏�5���tr=��L���z�_��l͉��dn룇�\��.���:<��<b{�?o� ̈́��m�|�h5�e�����V�E���e�/l�FK
��g.A�f�?�\<�����PJP��!iܮk�0��<��������/|wB��1\L[b��T���̃³�ʩ��ߜ�S!����tٶ�x�t~��rR��$�)�W���J�_�y-��9o��'�����+��UF!�O����hNݩD	R�ˍ����;\h���T�뻛��ɇ����3�� kJV���v���(�M0<q?�9Yo���=�� U����@�B��rj{�����ʁ����ڊ�TS��J�c�=��OY�|��@Nif�K����>	�U]ռ�� �K�������G �˼|zgWXF�Ew�q",�T��=M�����>���=�L��3����a
9���1du���`�%p_�m��}�G�-F�����1�@+]�P䋪���g^��ԭ��n\�����B�m��R1\S��TX��>Q�1����w�]<�@�؎C��/s��gX�V �
z��>�X�	���G�c�g8y��6e<|�
�9�U��wA} ��.-1
���#��e��~jf���ʚ��|�鬓��#(&4�-���HD�c+�p���� �A�
�����Zw� �UUݦ��!�r��տ��<���Wl}��e�����n����o*x,��D#�+�	;����K�n\ �VR@8@�&[�����<�zh��ty�O~d]�#Gϛ�K�Ay<����w'CZ8CC���1�Se��e"�)�śmC�o �5����fy��\���e�4���i.�7#��u*�����7�A��%8�c�df��n�Ư�C��9�< ߏ�� w�P��؁Y���֞��M�`X�'�-�����1�r��@�����TΫ]l�7`�D�x�Mq�A���w빱�m@E�><�`)}z�/=�tnSg=��@����J!xƧ%��Ҥ���x$t'[#�� c�!��)���m�`B7H�',[x~���iЯ�x��-���kA���l|�Θ+������<s��/v;�%L9%t`뉌8�����2;��#r~i�|"�}�ݎqL(s?[��[�ꮋq��G��የ8���jܳ��D΋��?^��M���
���8���t��������[;���?)�$l�+܎�	��W�Q���`<OK.��:_�����\�[���ۡ��є6Ua�c4� ���ܰ�?
T��ɎFi�q,��Z�����6��./�d��ŇV�/ �1	�����<�;��m�E<���\~�����E���t��&^;��u����Hc~�KnC2^���Y�w
⮒G�m��JB+f�9�I�cU�w�D���Q�ۜVV�_}).Ɗ|�g!�7@R_lDf�S���{����\{���{�݀!��ߞ�Y���߿Ȝ��U�b_>���t�X�`_��Q�=	�ݝ�˳C��<cE��X�����K��.�I!���V�.��(���Ȋ;���KSr��U̾�#��;p�A���4+R�we�|>tV7�Z9#B}2�U��յA����, ��6�`��;S��K�qs�^� ��O}�X��\�}X�J�R���	{������ZA��/7,�����[MM����Ν)Q��0� ����#e�?��7�z+C�'3���Z��wkCI�x��g��a���K�&|W@тG�e�+4�i���.�S��	Cڰ@��m1z�w0���)�+����ΐ��3J���|���RPz�A�ld忈B)#jכ
�c���pz�1G�{j�t�E�?/�.AH�ϯ;WO�GDꈆ#�)�N���N�#����*\s��
@�O�@#�" �a5/���4\�7��_EHs����%N�?�~{����e��*����Z�_(>Qu��벜�S��h7dY6��ܱ�R�r� �9
r)�\=��w��n4A@u!���{��Y>R�E$�����?�Fp�lu����ت~ U�/��l
��e���_dg{�{���>%ΙS��0�dEi�����a�:�����]��x��C���� c?|�|�)���������=�>������|�R���������O����j�e��C��E����~����L��u��롌�@�5]% K��4M�gz��Ht��
�pr><mT�����{��Nk�I�����z�/L�p6��ŵ���9z���:[d��E}|�D�.C�V`��XiH�CL�����J�h�`UQ�������j�=K��S��g�8�٢��3��y�=Xs�=�WOp���K�Ƌ|J�Ug@�=����1��P@Zj���?��Ƥ���ES�����f(j��"����tsVih:l'S�G��{X4[�O���8/�*���ң>�A�ψW���â.H��n�of�Ɉ�I���zVu���|)Xj't�c9��DKf]�ϖ���3��N�V���8�|o���������盜MkX/ch6f�G���)���Ĵ$=��f���@F�� @ͻ5{vh��!K��*1����*�]�;Ѹ�&w�BD/�����`�_E����B����R�2G��/ѥ&��<�S���o���%��7j(K<,����	�8z}|A��Q�������[��eNKq4����ip��Rc� 4	��S��m�=��"og��]��=�c��&'tf[68zR���5�/�*>���1�>(�?L�C.EH��M�)y����v��{��F�_�^�9R��=�r����d�G���h#b�71�9�N�➁��^ê�����~3����QIf��Eٛ�+�`��z,��-�٪��'QX(�P��}:��=!ћ8������]5���72���@��fBx3��q����M�3�E1�mRQb��؜Dݼ��`�Ӎ����Rڃ��~�Xl������2���^�Ƀ��|��������^��\�"��"�v���ٻd�Q��`��8�����R�5���ŭ�?P��'��KQ!{gX��Gx~g;��c�d֌�(c�0 �J����Q�u!)	��̘��#H��Z���$
�[�E����xU��r!f���2K����T�K ����v�3��J9O��R�Y� w�S���9�	�ݩ�x³�/ܟ9F�#��XIZ��ѧŎ���I󙿆�v]��[j\���pN���G��mx2�x*�n[g�Kc�A@��f���ņބ��\�1U��>Q��bP�7 C�I>��[��/���6n�_(MH�1u´�E���Fk�Tˬ~��>Yz�8y������V� .����3����4�V��p�T��:y���a�N��7-MΚ0K)��'.��Z��->��g��$��L����VϷ(����O%�%Х��\����r�������}_��8R�n�$�ء�*<�s#���(j�'�O�d%U�c+�����)���u'�I�t_�i���Ā��j'L6�V5R��3�m���8��� ⽩�t,���Y��{[}=�e^��L����f�	"�6��4��O���ɮ��QN��\�k��E�e���2^}��k�\�&=��*��������tQ�f�q�/���1�dd��K�|�$v;���S�t����������JA�X�wzH�����-������	7$:rM��rlGi[��t�/WQ0�U��*�?v�]h,R�ݫ��t���N}���,�?	oy��^Yez�V����	{��^�m�
��b����>�$tl{�u��-o�w���u��?�pf�a��4��5lۋ����6�����sܖ�z&���;ذZ;[
m���P��������T{���@�jC!�7\��f�!h�jϧ����xx����$5.�d�:g)����6��JsZ�>��ݬ����Rs�d�3����0!���7��	ѓb|��LRS{�o?7<��"��2V^x�u�˚�c&�G\��Z�d��
8��p�g���hM����6�8O���N]�j�Q�3�r�M9H����j��*K]DQ�����"��V�xK֭�?����v�>X4`�ҽ��,�vYn���L��M�.n��)�_`�~d�����qZK��A|`F}��`�v,}q���U(��@�M$K�� �Ui������Ćk]�0��(�^���]��+l�Q�������#��ԠV�ѡ!��ӂ*�b�V۱=@]i0�I�֙��و��[P}|�;�k^ ډbbe%B�L!}'u�ݾ������e&N���\̰14���-9?6 �M��C2����\�)`�o(@#sab)�@�⚁^�����Y_u/�I��Ȍ�	WɎw�Ip�tyZ�	L!e�KV�-���>iw���o�{ْ��I+��k}�TQ��mu�N�6ŀ�5e4`����[��Iy��~��3��K�ʹ��#�?mb���T&ѱ�e�u;�>��x�9&k�6o{� �$���ۡ������f5�=�k��z�f2fn�!��ڹF'�(�a���5�S�0	�EA
��TW�P��I�j�n&=��M^�z
��r�g��w���O���- �\dX��b@t/E�� ������*N�� ��<��Y�S}.k�>�Y�"4x���N�Y��&�c�����g|��r��ʽ�t)�}%~�T��E��	S������F}�S��Wd�����5PV2���7a��_9Y/��?�#�8Y����N?�jZs�6;�0�*�5��_넽ob�\`��zԟm�����~O�6�h�Lw��(���9�N<IF4\���<�M�,������`�{XCI���v0��o2���v�������x�	+I���g��jXP��FGmI�W���Y��J�H�S�"����;i�"I�-����,ϝ1�� a],8��"��!���kf���L�i�a�rw��~��?�?L]XT]�>��'���Āt� �#�Rҝ*��)R��1")�tC��p���������Yk��~׻��{�y��t݇�t�yZ,oUYI��p����v�ܗ����Wz,=l:�ØN�F��!����o���׬/(��2*iݯhyG�J�\c�U!�����Ub��=���������G&zФ7�Us#㗿[EUWu3�n����O�J{t0�^ -�џóu�0�H�ї�cl)��7`8���Y����y��S���s:��ə���V*?��d�%�g������+Z+	�P"x��V�g�)>�RL�΢l�V���s�2&������>�Ƞ'�.�����W�<�OI�8�f�E_O�0�?	u?YiѧQOj�ч.�żN�V�U�{44��9����^Ш;�z�(٢5"�x��1_�Nw�*n��=�L�iڼ����t�H�B?���4׹V��;Ԡ=�J�J	_]�n+����s��5K�~,"��>�=L�M�F?ӁV�[�uN�&��󢬨>�;<}o�;�aCc{�zf���E{wĕצ�%[L
�lERC�5Y�{�)[�'W�xN!��=MI���q����`�-_4[�f�'dCvc/�*{�z�;��v�ɏ��H���+I�X��TЋ'�-��sT��9�����O�B��^e<�j�gD> �C*'�2�7q=��H��^��{uJzQ�e澴A����9$��"���ܑ���k�����Gk*%��]���{|Y��!��Wt�xX����v!-��p�����7������}N�eE�̊y�}֜Fْ��k?*b8��!�L?��[�軛F^�j���}	��T��5��稍�_'�d����*�V+_Kf~��:l��!o�{�4ҿ@|(T�gU��'�=Y�i��L
<�"e
x�~��<�d�*��~+�X�x�2'oR�c�w��l���ty��~l�-�q�jq���TI����zӦU�46-BW�C�L6�� h|d�x���f�\�nG�#A���ҜM	Z�ٻ*�p��}�Ic���`�*R'��d������w˖nL��ic������o�6�"��ǥ���<SD^zB��{�ڠ�?��U�>�����l1l�A2�������O@t
1���BӁ�)nyxP�պx�`�ٸ`��xAQ�sJ�ϝ^��߰+��087�)ea2c���W������F��yX��o�\$E1H)6Һ]W��sȠ���S�����}���ც��D�\��1�&wy7�����%H�>p�劓s���x��p]��$��MT�w�]IPa���E]w'#ɓ8k+S��?������7Dٖ{����`�d� C�8�����^���aå�PJ��/iMnWV���^�Zrґ�H�in�e7C�c&T���f�a��PHP	J�^�,M/��ڨ��0;N/�^��Ѭx���<U���v���3�9��[��Z���'�a^�������~o~#c��-ȱ�S�D�f"FR�6�g���㦊���<�e%��YeV���J>@�	��QE��P��ה��4��%�L~�{v�S+��^�t�����[؎0�����O�齲@o�����WO[��~kw�h���s
��2C4����b�>k��W	�=��:�&����u�s=`�q�n4x��n����]��vi���2�雥�};�'L�{�sҬ;�r/-��H�W/�XH�|>��Ƃ1�� o��`?�k��a��F>C��4ǌ.ŭ��v���[�P%���H���Y�w+�"l"ez��l�0�H�?O�ͰD�~5C�k%�|�xj�W�iW�����=���5��<�A��l9�P������@�P��{0������Z�,�u16j)�T�T��WNH;%��'�0؊�d��@g��
?�R�I��w��ܡ�^�Z��@�Z|k{���Ѥ�g"J�&�ȸ��@���.�����W�l��yT}�?3���Ǽ)| �LW�.�RG��-��T]�	Hf�/|� ~a`���<�)W�e|�v80�1�]��鿰6Qhu��)�Sa��1��Z�\�l}k)�<Z.nmX�bϱ+�R���z�2��!#�3��Y��7���Q,g��ZA�UEL��ːG+��\�AN���pS��ӹ��fYG���o	V6�e��Ӑ�b�V��^s�q�1���'=J�{��؛|�Qww�0�A�n0�"�<<J/��S-��Rh�k�M~ T�ԅ��;i�Sgwˢ齷�z:��E�c����	H���[wᘉԭ��@� ��5ћa�_d�uA�/l����yJ���|��j��$їxt}�}QY}j'�b7�\�_d�&��yR���%9u���ܯ�Ť`��6�A��K�*��C����`��+�l ��0�O�Ҍ��aA�o'	b`����qe�,���jC_tT��~��!��[�;g���f�T��#���nFΩ�4�knkq��Ӗ�N6Q�6sf�z�%И�����>��f(��˝e�i�b_%R��ɼ���p���,=��"�\�{9��\����3�̥R�U���򻞠� ��w�S�rC�d���,���*���U�f�X���`�q�3g��;�����j�_&'���������\�g۰�!��)3L����z~�%�˯ ��](���BѶ�R�ےF����A��ـfbl�.OL�u�:C���ף�����X>�Pk�}&C<�U�}�KT-�Е�:���w4�<�C�뢠2<v�<����@��m d�Ӣ���-��I�:H]ۂ�E�ì%��)������!$�j7�tOcS��ܾ~:e�����i�Nh��Ȅ�����oű�Ȫ�Ȅ������t"{���[���%&���p����3�c�凰��Pu0�f/O���L�0��	gm7��5����%�xk~.�d"x�c:�۝� �M��eJ�Ҷ<{^r��D�(�R˯M�ya�xH#�^hf�EJ��n���W�<�b�2�Z���</ߜuFV}j�@7���u�Gz���ݥ޸��H��ԫ<q,F��Fg�u����O��'���3���^dy'�z�pY(���W���
�)����V��,�3��������i��װ#�S�+���.�RU�n���v���}�?�A�32�R���'��0
�o���	,�W�
��ܤ>��h���\'�J4{Tf�ܡ�_-a��Z��(�mVVJ7�,>w�!�"$b/�ߕ	�m�ӌ��}�9�lp�;g�N�-����p!�N��:ң[���"]�
%�Ä������^I���s%�N��ճ>��y�ն�A�^�Y<*H(�E�9��d ñ%�E���dl�iq���=�݆O���_N�\GV	N�Txe��?���c����(��J���(D���i� �o!�bfq�534���̾��~���G��{՛�\-�~�7bi�gvE�g��6\4Y�h�6$���5����,�(�LU��"��l$4�?�� -;��B�&D��AIJq��.���jGlsWAN�8pg�K��~�����_�t_#�Ӥ&��qR���E�W:?�5⷟�-�lپ���& \ bV�\8�	^���DS�D-�N/z�5�  Z�k7�<�c�ծLF�n�]9&��L.?�a}z#)�4���Utc��ƙ�xj
�,�բ{�P��C��� 0���s~���h7����1f� ����ms��I� x�z�3�m]��e�[�ӐV-M�(���Hx5r�&B0���5��<M�*}GB/�%-S�^J�ʁn_�E�?�����T�p	p�6J�x�7�O� ��:�[b��G�Xh?�w+��e)�C#�������}}y�a"�<��Lf�^iI%�]���.,X������g����'.__�Z�R�
��P���HIXc��a��M��H@I�~��8�?�)>l'����B��^��q���f�(_i�u��w�Ns���ۙ��߽>�����TM4���ȇ 	�p h��?ݻ�����NX��[��G=X�Z׋!��c��k�Bm�&���Pxꃩ�'���u`E���j+\j�9�ʴ��k�����1\�]w�1��U��7ģ} |��1U��>�o��^�f��[X{���\_�z��㑡_�b�ڛ�v]��H�&{��E���r�r�S��>�����+V�����͜�d�K� ����z��O�&�%ߓ�Lq���pO��3h�J�5�^R�P�N��q���"T�8㙘��_��*Eipz!U��㦭��`�	`J�k���2��A��Mv�π�Ӥ�����l]U������PyQ���Ή�O�����Se�f17e��)�U�ذER�P�y���1�'�7�j8�DL2&%�x|uJ�AJ�_�N�l���_N��!:�b���^\���3?��7�}���b�t��ߴ 8�(���^H�q%b��U��Q��IV\�h���J[��s�O�3�1��X\wck���qtJ2���կQ����0�^�&�ج�c�t����C�8���>���պ��`�Q��k���ɀ�N��2��9o��8�k:=��ɹ��/[ΆC�N9�E��VF�y6l�n�`E���1r,B���$�i'KPaE�յ:;�Ӱ����f^������x�T�P��fa;W��pX�D!GK�1��#��,L&�w6DQ'�^�=@VU��rTL:5 ���Ήջ�� ���$'F�����B Yr瘎���%X3�mZ��У~��~��^����ZͲ�Y�Z��R[���jz���I�z����j�ȇ�����J�p"FY��=�/� ��=g����o�IL�J�K%.�n���É~To��w��K��[Y�ymF39���c��K#��9*a=���7�$�"S,�\i
$GzU&6]IB�����+�V?ی?s?��M Ҏ��;'�՘�b�F�ԡ8�4����廧��:F�p��ث�Ҏl0���V��i�켖����F/ދ��[�@rzܼ�Z���A
T��i�O�O{���91��������ҘD�n���&�Q�.�#z�䏈�P]i~ޔ'k�h0;Q��4���z��2��u�M��ni�	
`b(!󩚖���_���x��l'n��o��.�ll�N��=UW�����Z��s,�;%TQ`�F-8Qst��i�xY"l�/a�({fV���N#x�����B� �U���s�Kvc���*1Q�^ɥ�զ�6]Q��w4ť�C$y���8eq9m���:�	S���OQ`A�����#���,�&,-�cY�C�_4�O�~|��.K�f.�\rS�ח)�t��@a*��h����~�t�Ӈ���m3�?�BD5���-V0^����I�����<WJ���U3k	�8�^'�Q������'�u�o�o� ~}9�jmb�?T&M$vNm#�����<~���骼�U��6�w��ĳu�oo�qƩ���Wӛ�Z�&/q�~�����:�ٱT?ž�w[7��#w�ن�#��+��'��1�H#K�	i���Evj��D4G�Ԇ�8��/g�N����<��$�R�z���{V�W�[H0oگ@8�N�*���mQ��i?F��T `���� ��A�xC삫A�#7i��jۮw�"� �~#�[���wv@�8	�6mS���z^�T�ܱ����B���Olh؁��'����V�5��Z�M���i��x��랄]��f�+�k_"��- �S��z)���
bU1����`�-�#�	a�N�l�~)��r�j{���ӓ ��pIq��1�mAǂ�z7�pn�20I�i�j)A  �x�@�'�����Iv��|���%�$�og��i������Aj��v�9�_�z�9ʟ�9���=!�����⯇ ��#�����_�$A�g+�Đ�hT�ֹ�
'���G{!w�Z�i ���1r�"�qqg�}x�]�4�br��" n�h1>���!���7�,A����ɿ���;����H*3>�ĄQ����+�sKM��A���o?�y����_�F�v�����q�%��fhF�[�7�<Wr��zu�(���~&���m[��|A��(Q�+�@����
^Ӂ%=F�&��0��S��|� ���O3<��߼��X�ظ.'1����\��9-�r&�;\Gy�'�Wl�9f<��m�q�2٪�$��L�g��䕩��̮�-����"A��lnUSJ�g�2`��"=��(i��U|Xfs�i��wA��2��1�s~]b�={h�9�M�=ljԁy�w,�Ƞ�k�j�;���Ɋ�`A �Z���0�\��)7رl;a��*�\���s���0�B$`���}�g�16�R�t��ܨ2���C�ů���g)$�C_L��դ��wAE4�J�V�xڶx��
b癊���,�竩i�g�S�,G��wg��zq�R`^8�!�F����g����{��	F�R,,%Mm{AX2u/�a}����� �vp��XA�X�޻�8? N�kTؓ`ֳн�M�	�*�<�?�i?�����@�8oZUQ��p�H����`V0j:ާp�X�?�������P���W��`����}�c����$�	*}�i3�;��W��S�䳯��݃��d�ʴ{�[^�+!�A�!�u�Q}�L45bH�99�>�ɕd�	6��ٶ�-�T|l:�Qlq	L*S��ؾ����c�Va�����obw�H��{�s�{��Z�3�g`u2���ꙝi��_b�J��[��~1N}�W>#�Ѫ�3~ v��W;��ÇЂ`l�Sy�́�`s�Ig�d����˗2 �(�/�B�
���RD��ގпrd�MAR�P��"��%ﯔ?�z p�r�$�)��_?���]�`�È��^a�6ؚU��ZR]��H���v����(W!���l~���T��f_c�-F�Ak��K��������zn)���ɸ�}{9ixK�=`	��w4���23~������������|嶜�/��6�����Ua� ����dP_��"�Ӏ�����2������W����!���vnЂ���k4B�q#!�zJ��������� ����Y������8ki$��n�����MW���2�,���ˉ:�-1�������wH��Lhot"�F���~���/�5+!�N��+x95������~���Oz79F`ހ�F�\	좯F#��\ᯆG�vOTA���ӣ�@�4m��_e��\Z�;j+������f���������b��/�_/��O���9���p�?ɣ�ѺH���7;�hp����k��_{�>Y�d�������`��G�+ �h�w,F�����vX�n�+�O�>�����B������4;�'�2"�M 1A�bMHt�{��]���W��/!�?�4|��L�EA����H����GV��E���,��׌��7��t��|.oUSOз� ��T_�������ŀ_?�R& �}*�-��ʾ���{��o3��ͮw(��X<��_v��A~�Y���(��m�H�i޿M�'���C�����2S:r�$Ȧ%��n�C���9�c ��!���/M�@�;�mKtڄ	��X�¢7�@���È���l ���R�h�X��&@X�K���U��E����&0����L��3�T,'W���u�;�|vJr�ԣ���ku�j�7��(��)�B�n�O��J�J�����xr�y �F�$, �r�p��i��Ҩp�i�JW^#O:��流�=ы�K��,i.�-]#�"թ�e���W������xbn�����Ze\/�t�)�<TiL�V�l���](�T��0��"�x�š�<����RW�(p��0�3OL���E�]�ìx�m�$r�����_��^�5�hv�n]���P[�M�zM����0��S��N��G����m�%�SIX�=����R\�f;S}?*��4�;��:Oz���{�cٶcm�&lY҅K 0m}j;^6�[�_ ?�7�C�3U'�:H0�F�m�-@��72�CV�[�7����a��i_���(ү>�O�5�?��0#ݤ�pXL�i�����ЮoŤ7U���+�	V�j� �����I$�	����ɓ�����V�8�</vt�sd��bqB����%��RiN�re�6�q��(�u��S�SL&'��Ư
��1si�@"�U�&�_�C�XT��-�(7o>��� F��r1Z	��YD=O�F��b�*z� �2|�N�&�/L�}�3k��br���O��x�L�j[{3� ���|�=��vd�J��}�Ԙ;/>�kKڍ:�D�+.Y�isW����:#5i�2�D��XXI��K�Lh�rꡒ��* �(1�+�.��!���~zq�{����2���]� y\�ί}����8�]q����0F��/GQ������L�l��e4��ܹI
߬��LO�pޫ/�T�ӓh�K�UYb���T���	ar-ʓ��-|ɂ;�)����BH�~y[y�+��"{���5�,��Q��{s�ը�<��KO]�<�[�S��L/�g�[u���jNI}��B+a�%�c��FԀo��A~�2��p��e���~�t�{��_��ޜ5�����Ɛ�Ʈm��p�����G/��];�6}���V�q\ xD��JJ��u
i��|�i�X�8A�rL�pFf"d������I�P�Cj�u�vgh����y����A5
��M	,BXa�ǹQ2Xŕ�l؎�"S�\����d��%&^��R����WtO稉�+	r���O��T��p���`&@�ۡԼ��5�D�pN-eB`��&Z�%u;��U����Ŕ�0���[��+',�ߗXbuM?������^��z�_�b��R���as �V���Pc��BcQjd�ny{	��?��j3���W ��K�XǍC��ݦ%[Ը���v�7���K{�Ԗ�dl>�>$��A�lˑ:ѓt(!�_�8{a�g��xs}�!aŢ����2:HZ�������b�����U?���8~���5N�a�m��ƞ'���?��{�Z��a�O���fTX�-οB�lze�kW�����Z�d��k�r_��J����7�?������_-ay\�J���N�1>�1��!�!'�Fb

��m.b����?�:�W�q�V���'�s�bb�<������-��Ɣ��0�{`��;82S�~��ꗤm�������W�f ��$�<��!����#۸'��Cc^o<��_����TwP%�vWG�	�.1!�6�@#��;����X+ȳ����9�M�x��?D�G��o���dz̒i��MMdн�Y`�<�t���j~�U�n��T	�K3~œ��hUS�8�-T�^RxH#�=KVm�p2Z� ����]��qI��HSX�!��G��{�Jx
� ��>�q�&�����&;
" f-qs��`!~��|X	�c��n������'a��+Z��u�̫at<�cXrr�YB`W�zZ��	�6�]�y���E�e��LA.bN�!��� :�s��i(���%e]m�,fy㲤� ������~*^&��w��X��#Mω�qeD��^Q ���&��� ٨��%��Zu�K~~�h�m>U(��^r�H奜��Z�"ި��P�PP���/�d�?��N���Eª��B
�U���Y�w�z8�>�����i0MV�C�d���4�%���4�X�\�ػè0:nw�^�+�\X�e�EWņ�GD�0o:���7�-���֍xRGW��������~�z�hb�^��W%њ5c�	�I����~��9QwU0�{E�_�q ���z:}'-2h�ҝk���̱r����6�BFCYt<����Y_!;��"W-��yvw�_ȈC��RX��[���|*V+�9.ߦ�9K�u��֯����, �T�D�5(r �[���aò��du;�T��$ߞ,7��
�$V%�P"�\}f�s�����M
�?��:I�XF����T���`�|t�s�e�* �ȄP��<��8����&�sL����(�T|v)������q��u��{ڗ��
`�?DpxW��	���gn���\?hC8m*�t�!M�* 
e8���4ľ�2�\���>ա��O�~�럓��U����[�BL�#t� q�ܑb�ɕ�at�#=����͕-�Hd��/~�rh/R���� z��r����L�K����q��V��N�~+֐�'��VPSǛA��+�)�&�9�U��jo/��V���2�q�����Y�	��*�о�SEB��#%	���PcXn��]��k`B^$�4�U�l�VCi�k)�p�M���<���t��H���V������Tfkx~K�d?�����r�1���tc���F���l@�ۥ0��G�.�����6���F�N9XX�'�]F�����A��Q{�(XF��e�Z��J�;� ;��&)�[W~�����-�4x��#ҔƼڴ-��S!+4X��MK��yQK��=���<<�D��UC|����+� �O�5�E9~��2 uq��Or���r�ݪI���x9lC/9M)B���3g�۵/͟heF��%�L�0ul��
��O�Ը#�z��?�%͒��T�F��Y\4
}>���u�F��;5��a���Ϳ�䓱�����@����K?����7�� j�9XsL���=)7j�V�C����R�TKʸ�HC��*P�����5"|p�c/�κ����a,Q�f�u�y��ܺ�2���a���[�[Ɨ}��¾���[��c��K�xP�Գr�Y>R��0�zj���1�o3]�ҫ[��h���ʳ�q^q�f��48!0�̌��%��0�V,|�g0��FR��+���7�A(�:��Z�~�/�^�u�7��Ndm�7>��Z�Q�	��$�X��^B����]~���1�D�I20����n�i�����q_�n;.���`��Lsp2<?��?m6��_�@�,Y��xR�J
�`iFbp'��V�h��ï��e��џ�&%�Ь@ë*��@�`�/�5q!���q"��� ��ѱ�t���!q�/���b'��	"�m�h��N�{ ���nԪ��SV�y�6��`��U߭ۀT���Ah�1~P�S�RKAvs��V���!�߉7�%��a�Su!\[Q�f�ViI���4 �f�:5�r�I1X�7���X5�T��vKm�잌JX�@�{�����YSB�K9�&�f���r��w�<�K7ln�AR���8�����cƙ��<��/T����Y�V��V~�g��6�y�ȋ[3Ҿ�kuU�1a��n�����̖�r[	vX�1}�΍q'�?4��jC<iE㓪xt�02��;�[�өKt$��xR��^�pAQ�e|cK7
�����K����x�t�������${�f���E]����h���T0����k���YW��n��4@5'f�T1�I�m}=W�)j|��pAv�2q�s�N�����Y�u��#����Z�����C�l��R�?�٤ Xƥ�����F�f���r����]m�̤���݉��+�a�V�A:L���V�|ăy�ᖈl�*�^�_x�O�$��ޢo !A�`�	'd�CQOLM�1w��{P��ۉ��>*"����=Ax�Dr�M��}�8�h��+��^��mnگ��|�t�h4ή�
�������� e.�Q �$`��[<��e��v޿o[R�.�s��6iR�X���H|	�?wZ��U�d�+����o��M����Q<E��]]���ʿ,|�e��0�+��$6�Y��U�n@���a����@CG����α4`9��ţ��P1"lE�
���iyK j�}�5��|��d�]�G2�(/]����%���+��j�B���5���[<�r=�fB��Gs��BO�K�鉖@��,�iKn��{�Aie���
W����A�l�k��`��� , �c޳j	"`�Qx �/=�̫��1&���y��u>�����ci0��2�j��q�g��kݾ-Z����b���˓�������#���`'s�T�B5~��[�jC]��z��\�*�k�I�������i+�v�w<��	�;]U��v@��R�!�P��5�����C���eh�C5^�,.���^��K�Nf>c���L/�=h~��+�Dm������2�§�%�ɼp��ʓp�;�+ʓ��oi��\o�3/��tt�#��T�TBuLF��V9)�4	��9bX����62�9'7�Z��
|�t��R�Lm�#m�@�Y{���P�f����<�cXҭ��A�����-��r�xQ��0����-Ӟ@�7��,V�n*}^�k6��|�1����y��+Z^�qe=���k]�ӽ�w��?��m��u�F�gu�T�3�oN�O���y���	IaA,��+�i��BQ�ICE�C��cl[��ffH�3��kSt%a!Q�ԙ�G��F�{�)aKn�"�}!jr�[�D�yC�C�:ɤ_�W��R��y�33N	���:����ڍ��959�8m����a��������-���3�D��|-���'�sĕ�����헯����
;��9J����I�k�Hٿ8$���y�*¯@��Y�Z��b�]�L�<վ�����~E��MlR X�C�g�e��ﱣ��9�w^��R�����:�j=f�ms�X�J��%vJw�2�Х^�x��#>�T�����*��z�i�|{�Z�xZ'�a��j�T��n�؁y��I�b�4	`��n��!��Q�Ui��e�'j�:S��(^,��Vy�i�Zr�ڭ��6�@�1
%@�k�Z`�72i`�'���H~U_۔�>���%]�O*B-Z��_)�kXM`m��*Z*g�*���=�~2Y�g���PE���>�����n T����Y;���wM>�cE�x/��;|��s�F���5��Ϯ}v�f5�
t���ʦ�[�3,��K��f��]ف����bǾ�!�'f-l�p}�
4��⏋Zr���t�$m>����3� ��������x�J�\^2DAM�R������a6��A_����Y��Pf��oW�������,�~/�󤸯���	��U����܌�a�j�j�PS��Y��M��U��q�
��Bg
��arJ��w��Bvb�S�x��u-f���TUV{�H�b�2q�)텃���XBE�i�[2�L�����>�ʼvkǾd�E���0�>wN`�l�u�c��
]>?�|IZ��y7�}�#OϬ�R����*�����-3�����)�:St���N|f��a�G���lp2<ġ-+�)�[oM��>l�pkp�����곇z����-Z��u�g�]��-�rY)���e,Z*��(���-*Y��@���|�U��C��="�]:D�=K��O7Z�2���@>u�^MT|�vhs���
 0��]�}vy�/~	�^���X�mg~# ���U�)9y�eG�V�w3{fɅO6��SE����^$�xV��q�(V�;��w��6����52�0���Q���.5<�Ĝ�[�~����t�͘���lx�<s�d��*��ǭ�S=��j�w�@�5�a�9q��۽��!��5�����IA����bк��J��Ƒ1I�	��k��I�S�4rY�p�~�
�ë��|$��<��k#�3�������AQ���/G۬���d}T�j��ː��ZD_ty&{��,"e~��^Lf�\�\�$��|VYt�.�=�te��n���ʣ�Q��������羣��%��?��u�L��`c:��j]/�56�Y�|����1��������q��/��=-e�mS�K;_��/�u�9�c]�đc0}?p\���c(����8i��/�Dg�kK)|�ݭ`/9� v�e�Jǥ�+GC<�jn:�K'��r����a���|5����m�O�ۓ����-S�M��"%^�,OA�TJ�,N~J>�};Ov(����fe��K}���>(��mg5���^ q��m�	� �=��ql�J��u���̃�f޴&܊ʘd��3MZ��r5�ã�I��/=���wM� ���#kÒ���z7+(�q<��/��.y+�O���a��X�����Hz����4yJ�d�<<��^}�E�E�z��p�/�;��r�wI�����h̔l�(_�PVw~��a�/q�++5��X�OOG� ���VU�~o0�cz*�8��|5�s��3Z'�	�O�ۨ.G�Eu��NJ���P�`G)��us�����6�N��/d���I98����"���Y���ѶQû;���#C���[�7ބ�1�Ù#�"Bʈ�%k�g��a7n�|��?..	�������
}�4'q(�X��eH/���l��RǛ6/u�D6�QB ��9ad-!6i�s-2�jD�8Nb�}�Y��A�Z=p=!�M�;�I�!�4�VaJ���@3U:��t�9�+9��F���Z�SOaP ��]����BH�P�$�d�)��p�#���|{br�m�-m@U)+�=��WF;��J�_�MH+�����̐kƯ5T[���^B<�4��:�v9��u����Il��y,�
a�7�)�|7�c�
\?��9��@ឯ0Аh~c�^�l�����F	Tq�.���e�͓'��Ë0��䬰�������;*�W������U�3���2�EZ��ˣ>����*)��4�K\�.J
�'X]�ڕ��6��.�0�V�CR���z�c��:3�-���>����X�{���rH����;���q�pU��V���w�M��YG��ʦXl��9I�)��᫯h,�h��\w��h�h��:�a���G�g�Ki�F	[ʤmЈ����t5��~
P�;�_�����t��O$G��$��m�Hy1�Ź�W����Y4����9�C�ka6)	���y�?�QW���^7�f*b��&�������o�'$��"c��	�m��X���A5�J4�o6o<y��
:�D�?+�񉕬���(N���R���������މ2V0��o��u���ۺ�iH�漏u蓞����~O�ikJ��{�O�/�
w��E>����A�E8pMJ�z���P��+yS|ҧzv �*��&q
�(t��\��]�꼵�`�h��	8-<ҧ)"N��5z�������8�~��6�^谴q�Q<�������s^��m+2��*6�6�?>�u�r��Q��Ȅx����x�1$≵�JԚd��'���&}�"�f����i��P�t,�޽�xj�C;��63���"����Y��z=>���%ߣ2?C��%���'<�v'DDX��ϑ}|���i�����B�f��7�˶s×v�6J���"���N��ʍ�����NR�UJ;��9�T�<Kۘ���nj-d������!4�'Zf�����ff����!y_���?/����I��A��X�Ș���V�E����E�9سpN�c��w��V����r��-��Eu�=�/�n�LxW��i���x$��I���~&���������������f>�h�H����נ�� #7��#c��&�9g�v%Y*��I����1�BM`��[�l(
���ȹ�r�����v��h����.~��ܰ���nV�P[i$�3�'���HΆ�L%�ؼ��I/��Ί�.@����'�-�P��%=*�V��ޟ��BW���K-��G;0���)Y~[�0A���bjiƙ�=�^^~�[����8����7��o�G��
=�A��Z�LZ�(�Z��{�̱���&���� ʏ�A�M�ޙ�a�+(n����\�����O�u�n�a���*\�{唼�m޾f��g!�5L������p ���끕�Vc�_�����^��(V�a�����>�VަK���>��4�*�z��J�J��S�ԫ?��i��=�Y��FQ:���Ia�X�@r��� W�,���ޒ�e�]G�c��?��v���+���7�"��宽k�R��N�a\C_�&���fn��7o5����EVǴ��.����Gʱ�}ώ���Ǟ���� ޏ�]^�6�[��O��< 4,1Ie� �f�vc������s�b�\_�:�!G�we&��Ў[E�Cd�0a��Q���q������� ��j�C�}��w���d\���:�n;�5�fշ����CT{���/��%|9�w6��~��O�=����ώ�E0� 幏V��C�4l$�+��t���jw�8�ϧȾ~4s�N�w�����{����Qyo��F�]_In�j�;�E�o�ǚ�Q��:���=��+�iv+�J�1t򧭛�OF=�^37Td�-��"�N9W�DD<>��l77&8y���������� fB��1z��Q�������ȶ:��L[�����"@����Q���U��FA>��N+S���p�lm�̏������)��r�ޠ!����~9D����xJ�$l6�ʡZ�Ъ_e$���� *ٴY�(�h���L�5V�$�{���u�Lia��v���Ȯ�R�"N�r��x�ѯBwҴ��9�y�]�>�Nu]nc3���o�o���X}��L���q-4�߼cq��5�6w�&��}��r�[0l_�t�~�+�@�����M��u>�s}�m��e�ÿ�<at37_���J�f��w�#G��1�sD���F(�=��z� 97��.wL�3��Sr��AT!j޴�g�Q�kC�9�g���<r��a+���-�����_�D>���oD7~�����'���z\�����&�teWo�T���*� -r�0bꕘ^"��SykѺ�A�+$֫����l�;8;�d�P���<p���h�m�M�?�pd!�&����X�Cv�#)+,B&�S����dtٶ��R�}V^���α�X&}�l{T�|�aO�ι�ȈW����JeZ�c��y�it��}�Na��~oh�_/+F���a�]�dr�:�7�{#%�U�A5�C�L������0�PQF[��  04� ����R(��H#�ݍ���(!)�0t� � =t��5�����ޛ��������������Ϙ��؀�c0�ԧ�}�^^���$����"T2��m2f~��e/>���6�;i���"��#ۃ�f��#g�,7;�-? !�躗�u�=�߈�ܔn��o>"iO�抖� d��b6�/e**�J
�[�Sr�P�&����]Kr���i�d�O�y��>XM墨��#���}��b.�0H8�\UE'%5:���|��~��f�6�ڡ�]7Z���Z��F�a��O*�zL
�̳�7��mz�k�u�>9 �u�G@ö8هf�z��f��0�ʤ֕l�d\?����~xF�^(Ka�왊X�ݕկ�3���y�g}g��L�=u惿ت��:�pfĴa�Ed��}m����;���ԋ	��ݮ�
�sEo������'�W'��	_�潿6��o��q� -" ������*V�1L��� �y���嗇��Snt~\s���Kļ��~����li��,�3���z�wckYx�B�T��V���N�M��]|��CRa� �.Z�rR?&�\1��9WL��)�%�4׽o�䂸�[ۿ>��aNI��m�q9��pg���xV<�$������3Ii�+a��ed����?�6Mo�Й.���
DX�e����2�Dݝ�Y���,�1���)��Si@����sY���n����j��s)�_�|U=�J�sU>Q�6�8�-Ռ����/�Pq���ߣB#�p��f;?ҥ�J�l�4)q�V�8���z�g��eW�ȱ�Ûg��$W�C}{�<��.4
�ýYk)�T��ǂ`��,�qb��U�ڲ��5/�U��hu�b�\f��V!w��0�I���4 �O�Ç�B�bx����_�=�f9�y�Pt%�c��j�et���J�.p��Or=�jq�Z���,������+t��fa����N��ޡ�<�$�<ut�H�.��l���@nGw;L ��e��y�2��H���y֐����愔�T�����0/�?��I�a��Ԩ��=_) "�'�Clf#��6��a������!$���&�<m��J	*�G�т�CrR�A~f�է/[�ܻ;�2��ȟ����g|*r���X�0Ld��|�ٰ.yM-h��~���u�!@�~�ǜ_�>~Pr's[3퉖���Q�j�O
��3ˋ	j�*ic��T�s=�����q`�B$����DỘ򆴭�����':������8�.޹�/w��dn�9�A�8����CB�Z��Ti�kG��j��d�	��]^w|,"�K��;�?w#�:*�L9�r��GxRAI����-�I�' F����;�XQ��[��@�Ik�}�Z�Hp�0��3�� ������2���+4i��AA�� 2Hk�\,����7��9��h��kX^�GP�_��?����M�'��%�����,�W+\��n��.i���i�q�3���l������hW�E�n���ؒ���T��槰�:��FϘ�3^�1h囯����#�^�5�uњ��r)B#dn���ʜf䍝@	~��Ή�͕�@5�4�[��6$	/6�~T]b��l�bV ��5���k��#P���W�@�5�4QXyDɝ�C���Y^^Q�9E2��k)�;IR�nF��h"ۙ֫�� G�ю�<8r�M�Q��U5Ԋ��~c�_3t>S!��7�������3��T�f����JO_��R^��h���l�_�9NJ(��Q�a��\�B@��U�����Rk/�����}�[}�RS,m�/
\�������R�#�nV ۤ��q-�{S��`�;�6�"�iØ?�py�U�}
c"�ɾ!�+g�,�^� Wò�p.�&snaQ��/�@'" '�.�֯q\c�P��C������M.R6� 5�A$��7�T�S�!v8��C�6���C��Ez����0!ߧ �{ڐ5!�|Q���R�E�̂��+c�B`���W�!��b�G����@���,Rh�J�1��(��f?TT�[摒t}}��(��d���
nܳ��I1�R6��˨ڥ��	��rHs�O�i����p���@�r�� �Y�ye�b��Gg{�^<�����~�Sr�Db�	�p�S�� �c��:F}�k�2[6~��V����'�{#���)����Ug5!M]l�5�J�#J�UX7�m�뺔f�:�*�Fi:S78~m���5��n$k��$I`<w�ad	3`�d"�q�������$M��d��3y�u��di�C=5������L��3�'��/�W�ű�1�3^�{�ׯO�Rs����?�D47aS�CF�o]c�KU����7S�>�@b1���*Z�qh9����˰}���.�����6�!s�������X�{>�?Ee�w��.OW��<�S���`��X��:��q������ #+�O�������f������hxyw�֕�bj*��tSs���Ņ�(M	ڱ��
���n�z��E�_G���Q���CP��!�/��;!)	�����&��l�����Ղ:�,&�'�>i��3��Ѐ뚁ڼ˚�~�aey�{�^.H�}��r�K��vė�fnT�h!!5�D��/�W֝�~� ��#+�:�}�E��<Y���y�t=t�� e ���[g���|U%
=4M�OU�Ġ�1����L}H����oF?�NT)S��Lf�8<|랪qpCsM�o< v�Bsi�u2�3��p���5/E�4�&�	�9v��W�:����'�T����օ/�^�f���	V+���jZ��s���{Wa\�DR�$nˌ�w4���!Y��굧$��`o����Ă36�����\xpI�)�1OW�Q}����6n��������b������@���n�Ր~x�x1��d$0�#�j������*�Nؕ,�/˨ ��m�a����߁��
�Z�DŽ~L���Ǻ�e�7c��-�p�<4��i�<�	WA���`h�NWTۘ턆��n��dB	�! ��׌1��p�?�ffy�f��\V�	����p#0Z2,�ͧ����)�	��
�����ݙF+S��5��q��D��<��"����^�|��a���ތ�]�g
����h���[kN?[��"Pi, | TI�62Jϕ7�^��<��Jd,gY���0ɝ<?�&�pR�sA��VP0g�B@�8�Cgs�C�>����G��_=��n���_y�ا���V�yP/��VO������8sw<ZA��j:�iHo>� 3d����ȗn�QS ��֟��s���Y�i	v��р��P�DDx�Mh]������+��Ռ#�QOD�7f�rͷ<Ic��mN���y��Z�P�:����&w��̴����`��p�����җ���\8ۙ�1��7���n�J|���XC'�߂���s�mț�WGZ;��B���05*�C&�?:�F�&�e��b %��� �>�rq'.e�5;�ѡ9�,�Hk����jV�>�dٞ�ٽ�v=��W��gut���'w�9O��	?Bed�H��4>��	m�(K�vF7!cy@�F=��Pf�c�B���T؏?��r-y`g��:؏�qwn���G�A5_�~�{U��l�s˱⬝�C�/B֯��H�V�<8��QF!�����7�̓^À�zF(~��"�Le��"^��5��w���gJAg�3���+���j�]	�E�KpR���CO���f�	+�/uI(�Ρ]<sG��_L@j��2_��{^�EoM#oi���E|FH͝��*o�/'A&3F�����7�8Oy�&m�J�U�󏨀=У<���vqT�c�0�	�����s�E������:G�a��v{�.�õ-.9Cih@�m�8c:�{�~����Z�� �O_��N��9;
rԢ���ԕ�
ln5�#���&N��afWe��(͊i3����w˧��ժ���'>����{��[�kN�����X���˔I_��0�i��熰�<���g���ĉ�����I��b̪wr�訒Z0�H�Ϡ�GDu>��'�˙�f&y�A�l��5gQ��6�[�8 �r��_�\�r�Hh�vS�%���|�9Y I�B�=�����Ł�&�@L}.��d��Y,��)�iv�Wmz�ka��$O�� R8鋭��![-B !�!���v�]��Kww:���\���{0eE	�AM]����#,fzL�*tŕ#���)?��C��)z��d�W'+x:���`p*�	��*�H���U����n���m�����!�lĖh���Ԯ%`d ��^/Ai�s@���_*-���A9l78�Ù�L��>�̉�b ��低���|¹�f��'���hd�z�]�*n]��P�T�OB��P�_� ��(�=w����fcP��^�T~S{X�!��8��ۂ}9��R@}����_��D=hL���Oyٔ�k��6h���>�t�/���ڋ��^u�&φ�ڛ��CxqzyCӴ��߃ƙ��!iH�L�ι��gŵ��EN�R��hYd�Tx��L��m���[��b�+�4mJ{Z!�m[���0>F}/Iv� ����S6^��'4�ep밺Z��@ W����aý�g��Y$�+@c!%_��H�B"�ʩ���ΟunK���e�xoc������ڦ�8�vwB2ݏ�dM���C��g��8^�@�'�i�!����?I��%�U���<ٿ��D�p5~˟�G��CAHz��`�����
�L�Fs}�Qb=���b�2���3�S���e�&=T(��^0_�?�f�{���b˚�SwGîSO�mx#4oQ�긾R2��;��-��c�����)�6L�6G����:�/]W�	לz�3�3
-{�Z([kM-2Zv���x4�S�0`�7�`5�ˣ���`�	
��4#�`�����M�fW��4�Vf.�H�
��ǐ�\b�V���@Fh�({��ZL�u��JX���������-0���90<�8]w4��^fq�G��X�H%O>^�n�Fi��Z�����ۼ�{t]��ﻜ�0����J��&�b?�X���N���$!�=Ts�G��E�Ccqf�[�Z�D�DvƓ��gj̓F�w/�Y��Ա��\� ��c�g7ѿ0���j"�t��˕[��G�nU�!������"�F�?d�~X�f<}uVR'���Ʒ��o��:JI����5m8x�Cak@�P�#��-�öv	t�В�W�t�6>�c�R��{?=B7U��T��"F��`�����2j�i�Gv#�~��/����������^F2?'V�K�_�\OC���9�X��_9:�~�<�,�L�F��R<e�N8��W�1p$6)~��t�P��9����! :�E��lT5��_���=����BA��9�vx�7sV�nD8�%��#���[�E����}Cҏ��s�o�aLU~ @֍��6�7�H�����zJ�"�>t�V2�I"^�;���,F��O&�a��@?�����Jն2��*�S u4�Ak�Ո�7P��a�-�<N�Ņ���ʈ���P�����d� RQ&E���m7�ȧ�=�-O$e�IJ�uQ4��d-V�C7)�&�0�h���n%/�<������s2+v-2k��::��r'�ǒ|٦���t�L�->��������Y6nO��r/}f]H��˓V��1��|~/j�N ��{C9�3��d��E�߷o�����64byD��Fј�	D
t�#�ˣ�(F2�I6��%��9�$�?�䔞�93��4�O�Z�E�:n�&�NW�uQM߹0#V��_�s��Q��<��gه�{[W�&�\�g�T�z���&\��A�f9:���Izpc#���,X=�k������b��[>Yv�8x_-J#�! )?'��3c�f"�Ĝ �~�s�uuO?�6ܴLȨ~��wm��\�=�����k����1Uu𝹦Ēr��2�i��\"�g�+F�>�����U�M�&�����ʨ�����0VAW��%���Na,��S>��׿J/��ua��$����f�,�oy��|Ґ,���p���������X?z�e������q����0E�:�j)���K΁� `N��GE�P_}T������̩�L2���ٹ����zh�������K_���c���'H|k��{�<�>�ʣ��{������6j�B���+Nu��OZm
ѽ�zC�����sV����]��rمT�	��k���`a��o�4;�<�r\��m+�����1͖�a�=Pn���d'~C������g����Z<��ڃ%E#�φ\�3���b�{�G*b�&w�[�/)�(�C�M����~��I�3�g�60X[�Z�0a��E��zq�f�5ާ8n`�p�w���&0;^�Q��"�y��7�BpO�L��k%��;��Rl�$�MM�h�Y k�޹o@���Xæ�}�_1����|,�[��a��ѐ��w����b�{���/���U��4A��_ix6��/Z%ƨK�6�=!����[��)��(��c��<������O�-�3��u�w�;=W�#��TT�ۜl��]z:�7��rG�P�����f#��P����.Wt���^P�HH��)�tk�S}.�����
��t���d.]���,��w�����������NwO�lk�L�|�˙��%{�w�W�!]&t�y�
����rMগ��x�P��#W���D��"&o 0P]�bW�N'%�1��1�M	&��jrD�z�)3���T.��h�`�7���s<��S���"K�6Ű^�����~�g�pϛ��k�<�NX2Ĕ��ss��+¥�3�+�w�s������k�����̑O��˵�յ�ѣl�Q!s�s�����ɩA�L;O�$m�Qͭ�_�e�x���B	G�@�6O>����t��]Bj�ժ�NeB��H���oiuk�~��?�T�	��w�3v���6��`F}C^4cv7��0�s�/!�����Jo,Î4��\@����tĲ���z�
�+��)Ʋ�{	����}Ҁ�f_�
�Cܔ��R}cI4�*��s��dz�n��+�?<
OE��$~@"���:�Ǣ4J]��w�V�{�EuS�B����/ɸ%A�Q��DW�{�e!ٵ��s�%z`l�g:��1��>��'�Ǣ6��+M
u��=�#o Ǿ�@�)�tW<��uK��nS(��&��Rh�C�V�8a�ioR$�1@b�G���/�=|<nH��ԑkD�l0���41�'/v_[�A'�����
���	0��rW!�P���b\R,}��Uz�VgJ�p���'�܎��
g˲��[�	��]��T��~�3c��V*u�F�\�7�K5�G�U�c�A�U��%�0��b�ֈ���x�Ֆ�!٣ME�%��;o߃��6��ۑ Nތ�߂�X@qV��h��^
���r�<yF��
����^W!-��6�{�K��������vIX��J�IG��b��Z�������6H-��pK�Z�,��\�`�Sb[Ur�1Ćދ5�y{��
�����gE�@/�}��)<�ky�M�W�{�>2F�Ǹv��_��d�d��e�t�zN�U����@����*�]�V��۾1��k�&�T�����֖%�ws����gT�v_�ʪ��a���<��]�>OP����P�W�]o����~�c-��+�<�����ZW.qK��Ϧ��3�9Zm���p�����)[�&�8)b�OX6~k��{`?&���'E ��x)&��.�ĩt���ѭQ�Lއ�X
+��Uw7#/x����6M�n"2+�2m�:�$v4h!�n�}3zȱC��H+���9�_]s���ePHYV��Z�6�A���*��!.����v���1���?\�Z��l���:bn��5�H�H�X�wy�s��m �)�*��ް�Z��w�������Pj �U��_R��+2��x5dp���74^߱�_���îw�,�=�����0Ĉ�����hx�8�ɳ!n�Qcp�4$mA8*�)��Q��5;����s0H���Ҵ�z�����������Xw�E�&ɯ�U���p���cc�m���0"ƋQ�{P�Ʌ'�X�|d:����z4g�:�m����L.1F>��䙞i�=#o5�y��˜ٲ������Tg���+�u����f3���%'o��9�<�ó���O���a�t�I8��瞅)b�UAKσ��m؂��y�x��$W��J@<��M�$�sol��|�C�<�H��u�O+fa�z��?l<����X\=JZΙ��O�a�Ti���=FK�j��57�y&�k(�@x��G���l�;_����W՚�ۙi��:�K����?�$��"�_ZB�Q��	3s�	��8��#��m"�d�G@� �O��Q��1^�g�j�{��|�DU=��7T�#�`���#3���i��5�z�����y�f���R�8!S��ػ����e����6:�A�z��I�͟��`jǭ���_�'-H.���^�n9ڭy��-�o�ֽ.DR=����鴎f���-��#_B ��F4d�a�5+B���C��y��vi�;���s�r��d�ϛrP:��6`�����4j�'Ѕ�!��m�1��I_�Z%�~1�(�83������}��nݔ�Iw�ۉ
��2����>*���κB�j�*{��e�Mph��~Oe�.:���t�JP�圻��b��R�G1,g��)��N�މ��sg�s��sJ�֯9����� �1z�7��ؤf��AΦ��F����3��`2��	Ğ�;lT�N��n���쭭8<y��vB�E�,�3��-ß���w�e�ܸ�r!�N- ����NǺ<D�f�ТA;��*dt�zC��e��~��1�ìQ�VR���<���,�g��e��7��q��4����0�6z��J��Y���s��5S�J葻(�,��l[�"�Q�v9����S�}>� *l�g<1Ð��ɇ�L��E7�Qq^@0�lD��qJ|N���wU4y��;[�Ls�$���'j�Y�������{ҹDa��L���:�h�7{a6�P���W�|iy�e{&�g��w����4��7�>��,����,�}hyІ���_#}�^K��`�w����ku姃×W�s���ؤ�
��B��V\l��@a���]��M��q��$K�/��ݧ�ҷ(����+c@/͗���,��`�RY���D@���LX�K���U��+u�=7�8d��Bz0 z���_7�x�TT>�b��G����S3�f.��K#��������BD�-�s�z��@~m\�� ,d$f@/�Y`(/]�Fj)>:+�K4�i~�}^��*!�[#�]���
�Ȉ�� a�/����;d��#sv�rћ�(1��4(���j�̾�m��z+O� w��J�^u��$T:�	4�gnlFX��WoCq�������C�dg���$��E�}q���&;�΂߬�}T�.��;�{[��!�=! �5����&~/��{B�	�� ����Û��2+N�5}��AI9�#�o`�$P�6X^@#G�kMlJ� �K�ŔЈ��~1���zM#������$}�iZ�i��V�.�~Q�!A�SSI��Cك5.*����tp'F�Z�C�&K��936��1��hs��Ȍ.�C��X�E�U����s�K�#\I�bL���?���s͜@m]iO#�fWO�I�m�8�hIQ��]OH����.%C�/��1���:��5��Wfy8��s1��񩬈'�3�)�i����}����n�^ȡ�,������f1{��uM���9��rO�e�	'So�J**�n��$P���ȟ�}��ڂi 0�8j[�J�J[_��]��2�ڒf�.JS�(��͋����5��S�P�}�p�?f_�g��Vn0����Ŝ�d�玷3CЯ�*��s��#��Ż6��9�7���Pq�k�X/J��f�����R/���0���-������f
}4��m~z"�0���N�Bx�-5T�Cje$�ҫ�>#��Q�I���)<u�Ix���G���3�����,-��޽JG�xz�E���oz�	u&t^~o���B��t�����R*5o@�����v��L��8�����E�u)]���\S�,��qdUcA�g��Ƌ\J�O��5�rD8���xdL(�=��;vQ��`�E��w�L�����!b�E��aӆ2y;�WSʏ�j�+*�z�D��
�l�ߪ�#�*��+�ާ�~C��e2�U�?��Uz������E+7{v+��~7\��v�6���iBƦy8�]C�0����Z�Q��N��<C��TE7t��*��������	Y�W�낂Б�
�m���s���)G,S���*�λt36(���!lpw��J����F\�ΰ��ga�U�+ض�a�Zl9<��*��?�L�ҬP�~�v�͞xr Oy��G!j҆O���^�+Qo����w�^p����7q��h����y�"��:8^���r�(]��ŚbS9��(t�������L�	�;��*I_���r�}Ʌ�Wtg�6	8�@¦�'�8���A�P���?���?��J��@�W��h�i��!E{�?6��O��)�?��+x��1�<_�/#���/�z|��.o(�|c���k����CGpK�;+��ct��1��Ή3.���>��u�������Z�L�)�/V��؊��p�e�t-T�t��U�/���D�4l���'*r�w�R�~ ��] ��gh*Tm�R�趰����%���f�O�h~�%����������3@�DK��5����4P�?H�� ݖÅ,,/E����`����M�����E���AOtNc�\U�iۆ�\7�>�ZIH.���}:�"��+�M�vMH�O?ƦGu<+����*o��'U��S�5�U�ɑGQ13*���0����$U6����i�!�_¤���"1��8gLe��?%H�k�oϓf���[J|EY��D�7í
�16&�/�b�ٔ�۝�G�:�⨑��(w
�rx�3�3h<��ѹ��4�GU/����NR�Mr���a��'"*��p�.TI���_�3�Ħ^��_'q@�������zq8�B=����E�g"b�����b����I�y�s)�Y���a���t��H��A0j"[�������C�NG���<9��a��yͩ@��Om5�:1bK��D]��_���7W���~�,��ص�_U���͊�8�<[)p�5�����G�}`-�kP�1��C��W�y��PyV@\� q�WW���̷F�ɳ�@��Yr,�}��#'%����S�����
�,�n|�����<���h��@}7'J�$���j���l�����5��$q�K[oZ`��k�7�'e��S�n�]�aݘj�ę�k�آ�_	�y���̦�j���X⿿�}�^87�N7D��?�h�ç�m��#"\�ژB&K�6DMGd����ͨ�s���P_�k������-�%Nz˺�d�L���!����'�<��m%z�����#2�ӌ~GE)��n!.�,47�&�/L��q{�s��Ml���Xi�q�|(e�͢���/�`a�(T|c��?�x�C��2jؼ�iJ����G�wc�<y�Z͇�]�rL�/��Q1�6���O١�����d�E�1w�G;���ۦ;�������ۄ\|��WE�Q^5���T��d���ڴ�19e����Tb��,n!�7ӫ�w	�˽юӁ����-��#�����?;#2����X_�t��C���})lLo��_�Ȍt�ήϽ/�$=+ ��g�����Va�-h�k)��q��	�����d�E�.�&pm�i>��"m�r��� }��$�{�!`§�ɷ?�G���03ܬ�p�\���7�1ǿx�1�s ��s7�&��r�A¼;wPq9��i�S����t�$����Ɔ��,�G"���,�&�_|Z�6Q���6&E99q�l�-�Tw]EV��mk"�Թ�3	#D�홄>^={ S*D�������Xa�L.����\.n�]@Զ���&���w�mdy��E�m"��u]*����`?6̨M�������e�kN��]���H��q�m8CE��邑E�������}"��5�ן��M [���k�H�7sf4./���,̓Pq��e�+|����/���n�$'��;�ym߯�dB���#sx475x~�������k��?���b�8��b?�m�s�`�'���r��Y�wB�0	�)`Լ���&�%�ys�� ڒ�a�LE1�@�Ԃ��_%�ʔ��q؂�cg��tt9mQ���f����t��~�J�؀�
�4�,x1�Ҥ=��)�J�i#��� ����ͼ��Ѧ����D�f܉�>�N�	c'�D�%�S,��2sq�\��2�D��?�*���ˬĊ2�6�=��O~�n��ѹC�'���]F�)��a�5_pE��&��c�{���t
�ٴB�r�0��?��>�l�3��Y��ad��]��X>�S���O0�㧶:���2�'�_k�@��a����<#��svk�|�^4U��N�r��/n����B��$�W��$�\f��*�~�eh�:y��$[y;�L��;�~9��S����H`N<?������v	������L��ߚ6�Á�X�H]#��wZP���b��`:��L���c��ʟIJ/�@�!98�@�����2�4á':C��ӧӆ9��76RӫR�-�5��.��&���	�ž��ge[�}� ����߾�{�ZK�ul���S� Mu�����fU?g���iH )�X���ئ�C�i���D@K��G �\[����ܷ/|��)���A��TGVA�Ӂ?ԝ��+7ݾ�9��*=H��w)z��PN�������X�!��3�A�TeF'�;)98�麁f)���ҐCD��8@F�[!JS�K�<N�Ys��|��}�o��,jz���Mt�Y�&����"8���Q��-.����BEp#{����w��K�g�eq�}��`-��.�ל����w�����Q��BO6E��)14��S�(o{8ȰA��:>g�����D�� �7��/���oM�婎>��}��dO,���@�C�~n�C��8ww��,@&7n� \7��o{2 �p��%4�JF� ~��E�5�w���j�,�S��g�K������o����}�5��:
m"��M~,m"/�m���B���w�p��6}v<�_��Q�frLW`�3o�a�h�Q��ؠl���4_��}S�z��¼�D@���fĊ��C���\�ľ�}﹒{&��t�[l"%�����:�'�bB��}�v�[%>ﮌe������vA#�����$�i� ��:�r��܏<ɿ�fl�k%�@m|>R
�6J� ��5m�w4%F�^w
3�-�y��
��dc�B�.t��>l��h)�o�c$����q!���|8iVS҃�?�p@��M�v�[)�)��ReD�'95�uQ�<к.6��Y�Ǻd4`I��sJV��>�;�8��/h2*���脼�Y�=T�c��f�t�K�B���U4��-��H�D���K@���U�4¨q���pb
S�L����FgGA��[��d�XjW������N�������[ ��Y����#�p�2,�3gjN�kN<�������TK�v����T�{���х���gG��|� ����SE���'�߱Gft�+�+D;���i���u��-�?���xb�(;٬����=}�,��b|��|!��B�&�ˀ�A������^%m�L��I���V~Lu����dIH�8�F�JiZ�%�f&gM�1�w�.�"K�Q���o�JO��l��А�/Aʴ]��#%i�E���!K���LC�,���;\�p�i���]��� &q�P�
�?��j���P��w=�b�#�r�݌��B.<MS�ƽD����Ay���Z1����](氛У�C��3�c�뢯�m(���׶1Tg_iz�]���=3>�'X��0CD^������ �e��Ku2��h��0�`��|�T���J4*��4'���F�4��b*�=�`*�g�|�Ȩd��UG���͊�e$���7�{�{��fa*}�Ro�O�U0�op�`.C:�=���`j9���M��G�G���KS�Qͦ��K�
�Gί�����2��;�)��G�'�.p�Lrv��״��F)�ҿb�^qP#�J��r�� O��a;��ot�&�ӠA>�6$7�+������������({� ����B�⩓�o��+���4�꠽)W[D��i8�}�F��Z2܀l;�U�x���r���)$]�?�gV�$z�7<��i�5��!�\)E��~�E�� ��F!_����<�-�$��Z{�']���17Z�g7�.Tq�w��ƴ��غ���jU���9�K�5&/�0i #*�l_Dq�b��b3�ue���S�7��<�w'�������ǻ������M��2���@�?�R`l�=0�D���r�\���4.nJO��^��@ 	I��6�K�d��R^�dL���1d��
�p���~ޟѫ�'�2,��֡�n���nG�׭ޱh� ��헎�Gi�ܺ�l���m��YWL���H1��0C�a"�͕������o���6�����-�)�4�����>%]���ۂ=�:�f�-�ƻu��^��O�o��#�U�
?��Z����4���Kdb4k9ojm��_ Fu�~�ܚ�SE�=v�R�t/ԡQ�`^D���(�UQy�#�s�ٝ��.��x��Su˃g��V]�ɂ�'ڴ��8ˁh���RQd����c�z�BE�
C�鱯�M+�2M*�jf4(rِ�>
�}��s۹��41�6c֛��h����7��3�����dF�$�k��d�n��(��}�W����JC�:)�ӱq~��p��[�����]%c��$�B�����=��HV������{��,�nr�E䀘�4�(-Ot��}����O�C����!��?5�2�c��_fR�#�����-wU������Z�lvv�*��,)�6��%Oa.C}�t�ay;�ۓ����E��i���Y
5��냴�����-�f.���ԝ���z\~��s�
�#'��3�t7�_�8_������V��TKQ]U�囂���K�93�����M�X��?�m�����$oY�j`�O�&�qˑ�>W�^Z�϶P-K��]���-I8Q��#���H"H���h���������`�zM٧�Z��n2�fc�y�"�a�l�m��C3�P��'�ӯl�.d�U'�X�hߨ�4���g>�[x�.p��|M� W������9�s�ԸJ���3������!9�U�\��p��5�ā�D����\R&��=����0���1���g�
�r�o�9�����\�sV8�f�0��#��4ɶ`�amb8�1?��V=�,W��8)�����"�ل*�ȏ�1sB����6��fG���m����5�����`�,8��	�^n9Mzգ:�4G(����X�FE�6���U��3��v����^lb���jF(�&FcK���B����c�2&;�dBi~H��.v��f��׾�a�(H�^}AF]ۨt�k.�hڕ����Lf_;ck�A���dVl/{��[tx��h���<���Q�629B�J�a��V�v�
��=�QC ��v�)q�(�k�7��{E���*�4䒙={�8�m�_�H�@� T2��=,����/���L�7A�˲����Zp�:^V�8����?�S���*~j��|�ާ�[��uJ�sQ�ٹR]�w�g\��N�	������]V���t�>�q����юitм�N�����/lX=l5OZD�[PO��;��+^�@��T�G��K���=�X����x:MV���h�,��!�x�D�y~�����a1��f���$R�Ig�|��l<����suvD�C_�O�ev�ЩQg�^`w�k3|"k���Z��Ԍ�pq�4��PSӧv�%����/x�:t�%]V%���˙��>��b�� �S� ~d�i���J3���i��B�W�\=���z��8�TGI�s�1�����R�{���7�8�}���<9��V�ر��F��<1|E�({Bd� �k���Zh�f�s�u�h��C��>S��т^r$D��b�j,F��e:.:���V�i��1>Z�W�q}���=��}�9�.�<C�>�ޣw�U3%�X���ϣ��[�̺s���Ña�wI�<_�8�z:ч!��N,4x^G���T���.�m�d�n���b�����M���>��ݲ�7�t$�}�i��^#ƱG��̀�~��
����������L�H���C⒙z͞����c�����	=�9&�Â��ԇn���QuZ!�:����nE���Ճ��[+FTh'%��/��?Н�a��C��438�֘I�q�<����o��y-�v��,�͕�N�w�����x�1�P2�A8Q��g�^:����}r}83�]���n����x��mͭ��&k����=ֹqBW� ���n�P������vR����<CM����--3""��~��u�K^��i��_I�JI-���Z�4h��ώ���uU��\U������V�S �\[×OG����,1z���q�b��s����9	��[���eO�Un+L��r�d�\��bD��;�5�ܦzہ�܁��&𗮊��ؘ��6�
��c��z�����usԵr$CzԵz�yv�N�M����%���3����[xE����(�iP)i�a$	���ABZZ��K���c�A:g����~��o8g���X�5���y]�~��������ܶn\����c>�UN� ~I��9 'L���%�6B�?<#�8����0�?�)���g��O�id��J��_��x������n��&?��/�_���{q��g�|K���3�>�4�p?��T�Ҧo�]c��"��nE�|���@��ÝJ��|D���9��]#��l�5�݌(��/}�I2�U��\:�\>P��w��x�	�z�t��^4�y�s�^���z��gE�M�F�&o�@��/��{%���3dw ȍ�g�{��z:2(Y��h��-�p��5x�����Asz9
5.�G�����3U��f����@�.��P���r�a�iE�KMr?�ٽ�Q`�e4�������},V^�������E��/8#�h���Yiu� �y�m*����O��v�%�;��@�k�w%[�9��X��$I8ŘE�ORQ��� �7@)}k��~)���v�=���G���ũ8V�XF���6��SR(�c�����cc0�zmow��y�3�A_q���K&��L�u������u�j�)SB���޹��֮����zA+;���}JSh���Qv�:���F��!�?��5"�%f¨+���(�?<^�y�=Z����Zm�u9h��b�t\������7ҵ��K�͎ ���:��rX܄G	�x��X��_W�V�X�{~U��qc��lOO�y*I��d��������d7���;i|��P�֫�0d�HFwO]k1���徠>[�h��K���t���-oj(~t�{�_$�9��K�s��'J�W��D�V M-V.	���]��"$٣ �~ ��2�������n��w�A!�#�b�0�=��G�K�]t�H�#�UQ��\��ь"Wzl�Ą׋���GJie�kq+��4��.�\͍e�ݽ�f�  �/C�FF,x)�٣4E��8�_� �G��w|b�V�^�q&+`�>�*+�I��ވO/�l/5\55��l����#p�@��
*C%��.H�
��T��K�o�m�x4��L�!!!O�)�ˡ�<��%�yak��'��$s����
.�L����gR��y��h~ uQ�&��yF�����nc�s+E�}�������mgQ����%{�%�Ϻ����!T���6���N��.�=#5B-�O�2j Q3kz�Iqg���ػ7"�4Gvs�����I$�;�ch����.�4u���|/�k�
)��^���7������ ���3b�\�j�i���&e�	�sb ʦ�OY�S����d��l� ��t��|��y]��G�8����R���pl^Ǿ6�Q{����З�H�K�ВZ�r�C��"�����q��0u�]e+<��e���L��Q����k�W��R�J���)�=T1������x��R�F�va%� �W�����1Z�4w5�i��{������M+�A���i��*�C��R͛`�<��ez�4a�QVv��wW��޷Q��e�8�v�vk�C�ߙ�O�g��+1]�I��qc=�b{X�����/%���	��	r
yx�/�ګ����x���=W�[�ł�y��n'��w�Y}�q���r���l���������t��r`�Q�5���A<�7�$��^M�)�$	};�=2���6z��l�[d�_�n2���	Z���B���xY0�qG'C� �Y���Y�?6����N Yb5�'X,�v`LS�](���-��;H��Bq�ŀ�Mr=���{��3?d��p\��=���փs!LF8���/*�W����T$G:����E�9Kp�q�b45i{������7�9��6�{��estaC�JߑL���s���v5�u,���[ï�_���i�� $� gZ�)�j烥Q�x&{�6u�T��ڢ�"�.��%�l��<�1���A$���Ћ�~|ˏ����^��׎�����IBU!r�&��:��m����lGL|�T������?��G��m���*0�UW,�ƟX���-~9�2�)�N��K����j�����/���
�`�6 SDTY�\�#&YIm֌[�K{=Uc�,�"������?lޑ��&��w���-�cӉ~���n*�#'� eV�xK��v�%��%Ϸ1#���^W�~1�����5��p�=��/%�Yh����l$<����	EEP%���[�"��Ⱥ�)RҤv����~D^��ؖ���3�vW��y����`���nz6H�;w�Gg(�N7yy9�}ܽ��w�ъ;7�;(��� q��gM���Ζ��A/Ԃ�}�Ѭr��n}��sϺ򠏭���L������BVF�4���U6'��=5�">_Ӻ((�9����e�(0� dN�R������CyL�D��G7�����~<vDߙ�������>xd׶&%��-��mŰF7N�*|�sy�Jw���h�Y�I�:�MdJ8�����%�K9p�aC��LA�G�?-�T�$�׭TM4� �A�7��}�NP��
LB[�c^��=	s��E��cx�ʫ����m�3�J'7� �A]��`�k�%ݶ`�_}8�c$W�)w-�`����&��'z5�*#H7X9|����(9�8������=�x$�����2�2�~I�?ob�Ly��I���k%
�D?`{�<fx�IN=��b�@�=k�kp�ӗ�e5�ܺ��ʘ�&��O� A!8�S��1j�����J\��:l���	���p�����y��p�4��k��nl��[v���"��?%D����G�1���,1�"M�f�c�O��qy�T;8�� r�8.��rVڿ�:�C�#4�:�K��Ї��ew��;�hID��UM����*w�*k,dF9q�ߐ=X��][X'�n0��g$��$�CDMŭ�����5�O�*k��f-�g�s�F��B}���?g�����r�M{�W NBg�j�ͬ��f=J��@\��]\]jJ�Ka��T�WS]t�v�]��AS	����qA�\�� �'UDwH�C�R�t^=\�:@�X�ɿ�h�29�L�-9f���O���љ �3`��g����oq\���>�X�_e6�*T��X�mh߿�)˥:��0�j�cM|���w�D�HYjL�N�T6�4��A����3 �6��(y�ؾ��|4��T�v�[��S��f�,Lc'�݀��,MQCPr4t ��G��v��o�+P��˂��6&���Ԙ΀��D�_k�w��}�������<^k�9C8��In)=M��B�rC�m�	�3(u��5��}��!31����͎ي'�b�@�>���3�N1��x���8��tQ�C�� 	�R��]])}vD'���q���&P����-���5/�s���n2r�{�8��G[tqq/<,���L����|�	��.׈������[/�B�0u��M��#��2�=ً�����B�^?���bq4S�x*,�}C��k�Ct\׏��>
<z��}F��Y�M��%_Lfk�9�2�@��𔖰�� C����EJ���(�}��=�W��-���R��(���"(��DV'B���E�G�4�n��ɩr4@)l��%�V|;g��<ҘoW���pv��*�c���d��65�7	6ηW��"�W.;g�z��6Y ���O�MDO�f�ժ�{ �EE���������������rxgP������~f<D
�M2{�Xxm$6�a� Ƞ�i��}�7����fZ��:�触c��i�uϪ�P?�*�ڪM
�Ot�����ES��.	�A'��ϫ-I�A��^p�_r��%��[�-��ݯ��Ǔ��ٟ�Cý��o��)�#�m��+!�ӇP���_iu�����K�#S�8�t(���d��gY]��h�ʟ��]G��[���j;b���tW�kD�Z ��rz@�U o�l�Wt�쭭�N���;�;6Y����&��x�F��[�A��'�(2�73��"'����>Õ���8��Qō���y�P|����b,����^�:��V�K����L�R�����8Gyg6ֿ{\����km?	(�Y�i��'�����=��:��q�[>i�|(^q>[���7�����R�{��z�:��zd��u��g�Le"ӽR�z%Ծ��/�^x(���Ԩg���yzޫ��1qy@�|/ff�����s(�u>m5�7����sy�S������+���p2o��*�7)�����"ޚ�a�	�r�&6���_�
�6����/�2-�x�� �w�c��5�:���▉�&i��LJH�t�
��b��^q�W'����U�ã/���OH�为:�!!8e�=Q��pߴ�5�t�\PDG���xA�Y��?�N�U0\��-���sN�O���X�P�k����p��*�l�"Ώ'�~+�{���Qy!�-n�&�xCUz�WQ���TAd���W]Qdd�r�qn{�0vY�<e��mksH�!������a�&hj1Ur`�+$7�A����B���-t�P,�xQ�f���u� 4�,��>]@�a��k�o$�
PK�O*�K�ʬ��Q��ާ����_ceA�
�k9L��$��M⛶�)�y���=���Ɯ�bK��(�g���K�s��ޱ�Hn�+>���S�	!� �CPr��W�@90y���T��7�hX�r�/C<q9O���T׮��aN$��K�m#�_L�Y����]�F��6FjځB���d�u��	��)�j%��U^�*g��U��$��C�ܫdرR����ъI\��@�U��m���r�-��|��a��kO��ǡR���L���=�z5펜"�� ���b$��q��l�Cn��p��]��-�����Ea`��B�� �vP�#�¦�g7�/���T��q��1n�_j�@y�l����J�}2I(����o��~�8Ȥ�1�p�R�*����ub|Fl�0�
;濿s�k�+l������N��ʴg�]�4�!�dF������ͤ*�}O���>��4��������G�����5J���b`! �.>,��2����	�j{Dz*BH�>ho����G̙�m��ٽ����!Fٗ����3떆g%��L"��^ �oǻ��d�����+���n;�-��,>L	����l��uP��4�76i�O4������������Z{��{�R����ҹ����HxH���5Cv�HT;��|�oM�3�g9�,�V��4�U��|�9E#m��r��\��[}xQX����-H=8�ǧ3�����'��ԥ���9��z����K�O����V��9)<��]�@��6�<��c�l(@z��I��Q~o|��[կBI��[[�����I��}Q(�}�&�t��5��tk����O@��R��:,���iL����J�6�֡�!~�����gz!��K���R�0H0�%�g�i�8(uM������CS�C�o�D������P��9f������n�6De2�ϟ'ҷ�z8[��K�u���\/U�)�j8�Sn�ʟf찄��E]a~�.����M"7Cs��cC���?���L�2�J�� yR�D��H���l�צ�2��6�yg��g�>e��9^���wp%���U;U:�+Ny��K�v�/����t��k�+]�kt�ɺ�߻�~y�{��a���kzr�u�<?�w[�@U���嗛�k\��D�z�,fx@�G��H� \Q2�50J_�����*�����տԫ}+�4}�|�f�.��3O��yG7%Z@c����2���,.a�v�~9��~s���R�@��T�:9$;37���de�_\:zU��<2$TdܲB,f����o�Gi��n��gy�%a�`2��U,x��	t�:���!>Lp;�$S��W�6S5}_z?9�ϒ�sH��N��TՇ:���M3����z�x6�H�1��[P"�_�>]{��ǽ�Cl���O����h����3Vq�l��32w&�V��g�r�փ�k�����_���J^�l�����8�i�=�4�D�O�4�j;8X7�{;����](��o�@bn�ҊZGK���!��C�X���G`���>U}*��)�;�A8(V� ^�<mŸTq~��^�b�)3� ��%t��4(��0�s�<�0C� ��Eo��Z�pą���r�SÍ��y@U����RxF���JU0� �����V=1&���K3��@??����A�l��m�cO�+���X����
����m�=�.%�ad:Sd����������S�r7��w�.�Pk�Ջ��Oz6�Y�jz�ve�o�@��8��ɋ�L�Y��4D�m7 &����"Sؓ#�����f/BV��vU��Qeӗ9�5]�.��7\IVU�f��I�?`�uё/2�Կc���'O��@O��с��*0v�&�����hmP's�=MsKAM�Տ��Ki���}27�3z�Z��Jtw�� ������_^�o�J��}�\;�RJ�w�#��9IS������&��\�胱hM�&� z�W���>7���i�`���1#D_jUX�bd�@FS+�u����S�b�\�i��p8@��p���"(����F���twOl�l�Ǣ�W>�{7�,����dV���t��M���:ZF�WZ��f�J*���K~o�>�)+���=��3��`�펪Ǆl �B� f@@�q�Þ�����&������\���U̝�M� Sd7s�D�,ܒ���
���}L���P�Q}��M��Q����ڼ�~��4�Ʋ�_�"���}�c*��1QFv|b���Ύ<���z/��Q<��+犕��?Ǖ�	�A��9<�M>�T��^-�c�>Z�j�\�`��vӊ��1�����jߧ�U��N9�{�ߓU�2��a�ک���{6�7�h��~y���#H��Z��t~&�4]�r�a�TI���9�	�y�!S�����q����G������FRōuG�K��ro[�?�~L�_�A��`���nn����4?]���)߲� ��Ez���C��k�ϣ{�\�7�>����ƴ���G��=j�m��'�˺��V�㋕�&etvX �$�ͩ(�k�Aa�vMA^�Ί0?W(�� k�gӝ�.k��Z/Nc0��z/6�DҍT��H7Xޭ���Ѵ�ʫg�P�l�mr�gHS&9�GN�v2P��07̷G�2�}V����p /I����0� ��NW��1��Wg����w�s��1���;�����"-ܖ�����"DS!�Ov��ͺ>s�Nn�eLTa;-^��/����?x�H������颰M{%Z��Zδ�S�Ϋ�!ϩ����8iu⩷T+DK���(������ƞg��a�q=�I�����a���I25?��ׁ�F���:-\��+��:�3~\^�>'#��P @�����Ki\�je�j{z����H�����{�*�Z݋���rh�Z���°9����Q�w_W&2��-a��4����%Gۥ����y	���kHk��:۰99��+�|ը�c�0w�J�Y�4�}�f�%�[i>�J���xޥ-W�d���_��:E���,�h�T�+���ߢCԋciBf������M�7�pM�]��;��{��P��M%m���r!+�����S�-QX�*+��W��"=��i̋�2��]z���Յcw�R�,��_����ٻ� ���#�X��Ub����v%��}"���ȵ#�uj��Q֎�ל�*A$��Ff�����_�9%��:۱��R4��)>���7X��_�}i"�U��	?�=L��|5�÷�<m�g����>QB��y�g~�t����Z�p�\�%��6�wд��$,��A{��V~��N�/@��ƭ��Γ�@��4c�,oȚNM�����t����8D)���G���eK+ �MX�7�?T���Sb��z8�e̼C�^6%u��$ȍD{�}�~���B
r�L�0�]�K6��o�熵��>a�J�.W)�T���Ǥ��	��A�-�g#�0S�ae�i��૎�@�fe��M1-�^���8Q���Y�E������"��9���;i�gBp�A�d��Ҳf���FK����s���EMֹˉ�<#7<[� ����Ō��z2Wz1�w��2�� �Ѓ�������f-���\��`�,ωT�ـ$_"�]�1α����g@��ZdͰ�gc���+0�J���"�� .�h�@zztk������Q'�k �y����4	��ŏ�Y�㞼O�x�ו��1S( b��a|
Ϥc*21WJ�0*��6"� a�v�F˽Ya���P�/��z�M�GD~����$/W��
�V�?�k>��-80�v�F����M�)['���=�6jeCn�Ԉh؍ʀ?4��=ceq�y�}��1w2*��1�������W�$W�
��VJ�7���5���_��G[j#�(9}.Ք�?��yTh�2,�~r�C���]߳�(Ub%�s�s�~~�Nr�� ���Dn"Md��Ci�,�U}�|���2SR�����0l��0`�u=�U�7�e0����l8�ɝm���=+�dE������l�c��G2�;�&f-���.:����}~W����\�m�}=�'x�R^	a��US���3�@{�y�s�p��p|}?v�WG�������A'ܨ��y�H�����5xi�nq�����:��#a��*�+�������v߷�yʺp��Z���?��b�������$���3�r���L���O�-)�^�:0����7hGL O,	��t�X�G�ڵ���s5�C3�c�C��_�Y�q�v%� ��a�*��_Q���हX�ڎ��ӻ"��7���G��	�����nπ���69�=�d�O+�<w)��s��x�~�3)�z0���\��9?���S��x�$�|�@�8��V!��Y����y@?zr�I��,\�~�{*_�l�y��bEy�D�U�w�_��^\���7\�96n�Ω��Gi]e���H�h��ۂNn��>N������v
"�9��U�.���+�5Rr�8�0�������֪�O�gݰ�����h�`د�p�_�ke��3�$����EX�>F�&�6]���p@ۧW�]� �E���t�b������հ���h�r陉�<1_��:s�H�x��i�U'�g�l�����/=��=�5yX|�ȭ0%�Z8�q��h��BG~���[j2�mt�e V�,uԻz~*9� �m���Wͩ=~�hz�?�kq�m�{o�- �=Fk!����H�z�+��� E�t#}�×0���^��?TU��g�@��bC9Gw��F}	f���T#xg��~X����V�W�UU�'o���ZǬ8ֲ��s�T���yjQv�9s�2~{t�E�)��{Wbg�G��f������JT�|e�E�l�~���In�U� =b�Z��0��M7类���gs��!�h�yL5 a=[����G+�N��K�KuJL�	����T���{�F�����l���5_�yAO~��"�Aƅ�b�8=���ت���r����L/���MLn~�nF�Ib�g|��U�Q����U_��Ӣ��'�B�u�K�� "�������u�K������*t���[;�`�D����ſ�<���ik�<PmS�)h*�Q��$�O.����7�&pHTs,�>���L{ Oش��z������:1�%����OgVd:K衑�h{���\3�7��Lӿ����~��Кo����u3�ry��;�����켆�1D�̶[�m1@����o����-�����k&Z���olE^$�o�{K< �Q���X#i��d����~���>	�R�x]�}v���f^��қ�#Cr��Xդ��[^�r����B�������u���.J裷�k�m�{Z<���?�Y-��%�Ģ�@��nP��C'��s7=CmN/}/皴][�r�;�üx�y�qn9����"Z)��g�x��E|κ��rxJ�%P��[$[W�B�/c�/��C�a�q�ҧ��qh��]�[�"��~T����*%��e}�,/2,O������8Q�})�s)J$��	;o�l��ë�p{������4���,�̵���~��l��?OeKN��^�Q�hyƖ$�؎���ܝȅ=�X���0�p�=�&�J<�^\��hg��e?q
�;��C��l]��q#g�{b;�cIMKJ����M�X~_c�Zy����E� ��؂鰴D��┻bT-�bѫ!(�B����͑l��k��@Q��n"�WHO��_���'FD�W�+w�V�=���j����5�=���#"n���z9~�(��5AD���w�n�r֭��G��݇>�ku(���&(6gwv7s���s��T;�Pm;$��~z,x��r7:>P��Y��Zf�Ĉ���F����9�P����)�:���r�G:%�kf��T��	2��YxYu����#X�c��!3d-��s2ʪ��l*n���{�Q�6�ʗ)0����9�Μ,�y�x%�)T�HG�����a���J�z�_o3�h.g�� ����Z.��u8WtW�:,�Ã쳚��3�D愧)�6��ףy~cb��w���r�|z\zF�pkP2½��Si�	������a��"9q;:ʎ3����=�J��q��qI��]��|�N�J>rݳ��\�)ę����a)O�'��X���vU Yn�Q�~@���F�b��,n-��p���/j�)T���&�,Hb�}���	�n�:����i��ܕv�ò���>����W�iniV��9фy�Ogs���5	
r8���
 ����a��nS�O|���� ��}?��E
m0~����5���d��5�
;0�[)\\"���{�+�{t�@%9]��NiK�=�_,���\��D���`d����i��&��w��^�R�k��ѝS���~^'��SX�OTv��`���$��j~��M$m�0~U4j�`4�g�
�2sjd)�PU!!�HԾȅԜ�j.�P���[�ϳe͓�1�д���
�&³_f#*���03���J�r�t�hZ���q�I�J�S��'F��vYx5��6]�'����`��m�k��F�h:}�������&k��{��z��������Ь���ヸ�ca�;Yp����a|�,eo��r:"p=�~qF>![Ϸ�4�et3�!H���Q�h�f���cۢt�)R�c�K_�ݸ�TB��5B���yFlv����׭�䒶��#�����(}V�����USY js?6�^ C#��p�����a��ʧ9e���=	��j���T��Y���/&/b�U[�>ɽ�1퉟���_�^�:�����ye��Z{�� ��5ky5m�l����w'HC
a�k/��$����v{�.����<��T7ʞg0�Q�u�B��&�n�ӱ��Vc���]޿���Zy%U�����H�����O}���P��=����D5�r�hu=�!�R�7��}�д�D~�IjZ�A�P�h�r�y�x�8�9@�r��ܰ�h�a*N8
Yr�L��_*�9�]3r�0�$m���(���:]�Ғ�(��zĬ�y���g	>��2�8�n=��}p�N�B���m�.��b׮2��Q��3��� 9���Md�+@z<G���ľ���ͨ�`Z��6Z����������6JR���V?�g#!�����	��ص�|�c�jh_�%-��k���y:}�O���]&�!`D��;[��ZW{"P�,�6�+bR;7�J��T����2��?{Q�j���Ͽ�D3�+����"r�{`��k��2c	� ����
|�x;���4t���N�)HE���|w���ڪ�W��Ӧz����\��~�Ϸ��w��s0P�ٵ�O=�#��Zf���&���ͽ�&#��i,�p���s]M-⡕""&�K�X0MNn�dA^��]ʷA��%���^����,驽={���Wp��b;���Sw�яr�e��Xp�ܯ����ל�b$��u���=���K�$��u���=w�����,xsLa����b�s��V���*��>!�����rk����x;�$��~�f������)ȼ��t����2QX����(��H��SM���@�_)��s�&�|mk<i>xJ�h
]��y��c3&�]����AVZ��5&}8�6%�rV$�w֘�<���#�/3<��+������B�{�?P� �%�I�4�^���T#�{�&�r]�m�L�	���&���� }��(��h"+  � �ڮ>��J*M'���������h�5��^��x���㼥cUz�"z_�q�N}���Z������	)^aO� �$�] �s�����9�o�V�j��=!�u�n��,4�s*��f���/k.���E�x�~�y.c���R��l�%	���(ԋv�E�{y�3u-���v� ��j~��#x��Κgnr�"�@���7���z;�'���YX��?���q��(�����Ć8-��\� Z���w.@���L�hjҠI$�9�Z�>H&-���T�bN���!�i	V�4���vc��r���#�;���.�t�c�ܬu��z箯R�/�/���wN�E�{A&ӻ�2����m�tߎ���@2T0���ڶgE��l���,e*U�����"��LmU�qRi4&ą��3�f����{��9����!�B��ݱ5�+�HBa�%�YG,S���Q�a�>��w�&�h�ˀ�XK��;V7b���~/��亶0e�8��a��!��NB<K�?ѷn W��14\�]v�vV0���1d�NKT@Hf�ձ�*�:;ﭤ3��O�����O"+~�Ln�f"9�3_µ�&���%���x�c�Ys�VК�U�G�9��ɱ���ɷ�fۺ�4T��$�~6��'��N��v��~��5Q�_����J�|�WA|5���#s���>��̸��bl�Ϸ���M�sZFށ#}�9�P3���s�?����������� ��$�����4��0bu�jx���w]���4��{�� e�����"���
��j�-&�M�	�\=�Ͱ���<*Q�ߕ/H�8[�
QbV*��-\�w7 �^=��Ijl<��H��c4+Dn������P�]����{  p��~3���m�m�����D �KΣ48�<gA�=c(A�.D6��4��r� �1~�~�Y�|q�q���}=��'�R�G����b���[Y���&�����4�.+$)����]"4��W�>Z�{�.u�õ��r� ��i��S:{�ܞ�q�T�G�${c���$U2�8q�i����=Z���V��<��5/�&��M!^Ґ�?*��y���.���PJ�b>b��/\��כ���sOm� ��B����焾r�W���ݩ�b-�h޼�3۞�=%���mtG\n���x�d�ϋz�^��s�HP�C2A/r�\��[w
����$=a��j�����W=PC^�/)��D��vOD���j�t�<�3�S�OS�����j�)sf�b���:�e�:�����gm��aT:�]��"x7�9�3��d?�_�k=��b���B����l����"��~H�k@:�_���&zsf4$�"ES�k�x�*����6L@��o�
������/.]ey�7�o�*�=F9���
5����N��[���,Ń�vV<�̠�����l�4j�Z�aB=_8~�U��k��͛Ǔ�ʔE�җSZ ��9q����I7�����Q}ZM����ǇI��-5��:���Ȃ,6�a[w�0U*�np����v���:���m�j^����$��v�J�m���偾����ziC���5yeP�\1U�Jv;gfg�|����'iÄɍ{RB�SL�/�M@�(FS�ܟW#�q�9�ݎ��%a�w�n����W�Y���6���o��(g�7ۦ^oT%ǿi��|����ߡ��ҕb�wN��P�?�OU��j?ۚ/��q�f2��{˼����^m:���ǰ�:����@kt��a4x�P㿓q�e�c>f���d���)X���sh���`���Ul�����_���n��$?֐���s�0�eO�1��&lQ>�8�o����W�q�����~���fT����#յiG�i3S4�h���	���r�c0�~H�ؚ�>m��`ɨ�G���4*>#��	�W���_�'�#�X{;~�3�x2̧��ڊj��}s8闄R�F��߾�v����L]��tA�q����p�S���D"��=z[Js6��䱞���󥄭�����ͦk�Z�|e���=��{��r_[`�~Uߺ2.�(��eqd�˨5>���2�g���ɖB�~�5lO�pz!��ħW���G�句\��c���B���+����l,Q_3f!����jޅ\oa����\�w���8?p����,M�]�ֶ�U���T�M�N�9X����_��~�y�T)/���'��^U�7�q;7��gv�PX�ɆV�,�Њ4Պ��V,�k���(�Q����_k[�����v�'�+��"[��đw%39���@��o�&��t���~S��\�Ǉ�)Gc-�5���dh��dLQoG�e�d2T�41o}�v�웎�M������:g闿l�����=��c!$���R����=r�\i1�c��x��x_���;
q�S�B)�EJ�7����rP��}�w�Uݡ��KY^�j|��u�C=����]s�.c��� �|���\w�4�\h�',���;���p�ԓV̷l�ڢxQ��̎��N�O����>���>~y�K>�r$N1�{w�¤Sb������@�]��$��Es�V��ߨ,Pgx��C�}�R#:������(�ٴɣ��K��@��cq�����č�[ɿeu8i�yfC�6��I�<���K�.8+����)�3M%G�����{�4�g��fL�V�KOO/��y=�k�0zZ|�C��Xn��P9:�#0l����3C�h�������n��~?�|?���I<�Z�qr|T�̓y��E������������N�P�xQ�>S�)��h�s���a_���ƣ}�P�D��M���Y]ҍ}�ߺ楛$�U'��h��Q�wƠͯ�²ͩ,���O�ݒ�Ų�����%Y��� w	[����I��'N�#�m����_����ݛ''�A�(��u���G�CBi2(����:6��\�)
�m{w�6j���0y�C�����&����n^/�qK�uVV�3��b�䏴t��L 7 �*Uw'���X�����k�E����B���4m��X��ߔ�~�8h�+Ude�7�����Ő��S*��20ݤ����_?_�G����j�a�C��Ƿ�m|V$��5�s
�!ˤkl~qĭ�w��"v�8�IE�;������\���s�t��7Z��d�*"5c�k��Z�F��Y8=�g��R,�^����s#⛲}+���wg�S�_�K4:�s�ٛ���t��niD)GbZ��Z�w<���r���FA��S��ape�Y��>�DiC>�5�*{ja�/%�A�=�I��1w�i����,0&-����gu�/YpN�lG0W�}Y��a���n�Jw�<�s�d��5������s��'�z�����h�u#���������c48���;��N�1ݭ�� �_�vH�P�)�T��<K�̓��l3����%z�����rRPj���\�/�,1_��Ȫ�9����хӑm�X��;q}���֩�M/����<�����Zq-Ux�-ي���f��b���9;��l��L__��!��	��&ٗ�ꚁ�#�ܳ!�� {��@��,�"�n >&�&� 8��?���VեAf�벡���g��w\v�j�OJ�'��Jߍ�B�P��`�5�Xp]���%RȌ)�R�Z���_�ՔP���p��$<�1K�}�J�*����l6�:�3R����p,��oiS�I��&>��G�K��]�����,��Ie�5�/�	�u�P}p�
�w9�|�e�ڞ���=@B��E�F���x"̡~Gr=����NMph=ͨ���-���Ya��d��Ӻ�֡=�����[�
�!�����%��J�����Emˤ��.Tڋl'̵*�@-���ly�u�Jv��6�����h�= \�6�j¯u�y������]x5�6�#�g緹�����ެ�}§�&��^a��֔YO�C��?eA��c��K��OEFsG�p�V�ʳ��QGz��X_=
�ګ��'�7�}��:{�#X3��b�/r���&� ����?���NM?&���������k.���Qt�x ����Y�^��X��j�_'B?L�a�0��~�l�i�X��XF���E������= ^N�$K��������_<WX��;���;�QoI�agi��,�//�>���AL�i����6��W,�1 d�~3�G��䭞E�����q�0L$�f�]��랔x�ۓh���l/�W��lj����+�9Sz(��z������3�N�˷�͡�����fr�)��;g�����Ji0k��U��QG��9��O��&,�4��-�#}\���[{F���mi���fY��:.�W���*��AsΦpm��(���Y�/ot������J�;�!
$+U�(wa �0�`C*O����k����o$�l��[9)��gJ�����[�E��m�J*���J��H" %"���1tI��� ��RCwK����C73g~��9�p>�3���^�뾮���v
aV��x����U�g t⮎���0u�&5�~<:�Ysj���#L]���SfuK,�Tu��#���Mf����}?&�o2,rfp�������_I��xJ�@m���e�r�J��]KXj���b�Qӗ��x�P��B�̈���N�d�������w�����` s�6�q���G���A%���$��Xi��qL���}&�C��1���^�ɧ2�( 7؛qcu�@����$3h@�f�9��!j223����z�~@�M$���T�>$`���AF_:q�#��eˏ�W0)�Ѭ��f�P޴����T�H�%b'�c�$���g�>���Yye;p����b��q��1ȒTK�=Ϊ� �4��[0�m7���(�u��W&��z��3n
5��A�
�����8~��ym�?����z��!.=h�L�Ya|��M�b�	���Go}���@���2�/��\�_i�3i����Xl�{@���ׄ�/����hD�- q�6�߿/�3�kn$C�����U>��c�kh�Z�?��?�U��$'�kԌ⨝�9<�<�wKڵ��muOup3}3��D�U?J�F�H^\�-�7A7!��h��ߏ���?E�����W�yoW���7z�0���e�T�n�L[R�[}6O��C�ܖ�Ra�h������:Cw.H ݼ����%�ѵ^�L{��I���-)�Qw�.NHp��xu毇�QY��#��F*ۤ��r�[Ԏzz�q#Y�=�|�I�d�R�n���O&�jCp��mC g4E��4
<�4-��)�t;�/ψ�Q��˓����9��Q�"TP_FsA�xjr?9/����Nk��� ���d�0x��xLbـ~Ӗ���.'gz���pw�,�>��pp��s�u	7M�L�e:���!��+��ە�	@(<�1��vl~��-���f0	ͷ*@O�e+���NHK#>SAMHi3bX����PKŪH4kQ�89@�n���4��1D8<��z,3sA���פ&X�4��(���Hr�E�����N�w	 0������]�qƎ��z���_
Zz�f~�R_k7�oY=i�w�P��� �Ϲ�M��GlAS� s�X=�]�Z�ҧ'�mzT*/�.?��������=��胬�3�S�d���0����W���a���?NL�G������w�����E�gK��+\j��ҊzV���A�H���X��	�������l��0&b�D�+�Y��Zt�9+`�����������O��͒��Lu�dǞo�K0
�������s]�>rfLL�~.X�Ԙg ���]�,�7��&9c��7��Ă?^�*4�4Ei T��`I|���fcu+�`�@�T�G��P�N�p������6�Y�S�u�!u:��'�w*�3��t��mn�Y������jo:/�}v(���O��2T�xL�� ��h�
���x���cC�O&^y����ڈ��EN'*¿���=����b,bn�)��G��^�ܤ�ogѵ��������U3Q�����a��}�<�i-��k��'�� �����u~���ڛ� �iՊK�v��������r �v0�$Jf%>of@L�ȓ�6�����9�� ��R;�[�� �	���n=�{ L��@�j���\dN,���L�V_���}W���'vU[J0'q���G��Y-�)�/	w@�����u�[S]����Bu3�� oL��c��N�%U--d�맡�$p_�hl��kѬ]�DX8ϑ+����N0����pA~�d�2�Eo}+��Y�\��z��=�����7�K�UTQ����K�5a~�M�6���%�S�Ô5ic姱zAE�۾�ƿ��&
�1�%1�����,�7�R���W�b�c�&����K�DrwjkH��z�{������f�#��s�3z�\:��������&a37ƇպЦ����@~VO7BY�~�_w׏���Y -Y�g6�:ɨ;_%T!Ԣ0�u���F|�`
_KZ�U��X!���w��I���_٭��tO��E6:���O����qǛ�L���(��}�]�T������|���}�F�,�6c�K?D 2�Āj�yB�'�����w|�sw��c�Ӻt��U.A�8�Wqd5Q'|W�:���� |lu���1Z�ؘ�2�Xy���;�6NG���xNlE{jbǧ����[�Ol�L���9��P$͈\f�.����9ə��ot��"�W5Z%j�ً���B�!1�m�E��ǜ������7�J�Y�^�R9�=�Bܧ{^�5��F��O��Sl�[F���;�:��kQ����l�!i����t�4QoXo#���좩��:��]6n1]H�ۃ)�����r3u1F��U�/�Tي{��ܘ�:�*�:��K�=~�^P�3x}
�	�I��mt�f�CWHcM������QR�F�Píֶ �9+Mu��DSK��ߎ���P��i@M	����,�e�[��@�~������w�Y�������!��Q�|HN�yV�'����/�9�����u�^Eh�iC�J(d~��9I�q{���՞��i���65I�x�z
����pd+�Na�=��K�q@�E�hi���9jw�����ӫ�f 2�ܬR�Ki��O��soyA�d�/�/�e�L7�*a��=�$+f/�&�MA����hU�ߡ��_q+�̻��R�����p_�y�Q���l�ub�Wk��R�q��9�$ѳ��H�4�ʎ��o|��Q�$fc�%�	if�x�k�P��w%�x�[օż�:Kvd����90붬)���>�gWzܥ5��X�@��a̙���JIiӵ�]-�@�d�o�R	m�<����j]l����W+Ħ� ��J]x�A�E�SmL���C��:�gԚ��"?�Qg�4b��"�^��8o���0*���[:4N�ilm!@y�,J��}?q0�h !�~-��+�������p�_��K�q���:��� ק�^,�_��kQ�+�[�0/�T�	9P�~�����]].����	�F�H�C�ã��i���M�P�F����i��-B�!�]0����X�ܭ6��lt��Va�,��F�w%�Y��8�u1��!K���s})�L��^�D�^.8�q�Ħ?�l�����XXU�ySbva�����^�4M��������'#����t�J+8�*�D7d:U��U�~D����l�{�6�	*����զ x�?��k.�|�-���n��I�� s��}he=�c���D��>3�e-^�Þ��yu�vm�֣��l����l���n�g���B�`�3j8��d�gR��ȼ��$��?�ը�5�7{��S��k_W���(N��[D�<e�kGS�p�5�=2�Xo�@̵�}�>d��6�0��
�_?�
�Y�zd���m0�3.Nby�I/g�-N-�w(��j/=.�:�R�]��O+5J�[�:0�>�����CՎ���3�%N.���B�9��<i������s��c�M�z=L�ƴ�⏱��Ŀ:�+�9�/Nw��$�����(	�(0�:B��IA��%�]k��%S�D�'�L���Kg�|�9��j�@�׽֭��&ۻ��Z���xñ�4�ߘ�e�<>�9��=���v3J�q��\h��ȉջ�sG�`}֜�G?3I/;[_������SrVt�v��m��F�Y,W�O�@(*H���p_��.�֔i�#f���_�0���>	_<KeQzu�H΂
_����
��e�$�^o�A�9�6cxv�����v����ޢw�*[�_���oB=��Vc�Ǡ�Ƥ���ԣ\���]���^	>c�����9��7� ��޼����8\���Ⰸ+��DM6�'b�����UL`����^M@_�3�w3�tl���?W+������?Z	�@a'"!�az��s<�o\˄h���T�$������lGs箯�˜�Qw���a�oM�V'��$�>h�y�xx{��Y�� �@$��2q'�>�M�X>#6	
;D@BvX��CА4��y�<3u�M�@��S�&�\����������@O:v���^܈�u�w����X�B�ԤJ���Ʌ�Eu3ݷ�h�T2��V��j%�##� ��Ǵѭq�y~���`}����*M��I	����K��Db�_�>0#7Ei���?Ɠ��㛮g�)�vṘ������g���R��i�k�B����~���-*N�
g[K�K[D�Gp
���YZJ�6W�Gg�u�͊u��2�w�w
�B�u�� �.��=�M-i*�t�a�����#���u�݃�5ڭ�����U������rvR�W��eQ�������Y.bދ�=�.l'✁���Sg�OF��-l�z�ۮb�{�8C�~�������+���DT�%w��U%�24t����S��;�O��Ε�O%Q;s�q������h��򥑮yIt�0�U���{���I������X����)��2ک���&�A��Y@F�}h��>!�ԏ�O�9�>��f}�B:�B�q�j����C��� ͜�Q��<��/�D���|9��-L�\����!ۗ�vz^+���ʯ�Ae�ѐ���^N ����S�v�k���@�B<��Y���#z��?��BZe�Z������Zr�K�Gu��a>��n�A���v}AY9W�'sL�&j��e�.md1�hI��x������<��A,+_��[?�y�;��o>m�	�S���vz�F�T�q��3���k��i��q��FN�t�[�� l�c�c��6�FFb�Yv`�WP�����l10����/tJ����̆�g����jz�A/�+���q�~iXM&��^It�?}�Q�	�c�J-�����rW�e������&?���H�YF�3�ɚ?����wo���S*�.|��⡒PI`YϏ)f�8���}w��ҩ��=2}~�����0m�����0�����OS``7��_��?������i]�;B���Q68@��9E��!�Qo
�d�ϋ9�N#l��H�%�J6]�C�K�\�[(Iٰ�5��D�A#W��E�U_�(�ь�M�-�Е	�/�ٮ��FJ�j�(��j+Bw,��!|���}�T��dEy+T���d�>r��6�^�p(�ؽ�'Y��rp��$�8!�ǒz�E���L�V��h���e2�;T
v��$�=��;��<6��, 򛾬'�/n3z󗘁���@DS�lj�u��	��<�~ǣ_�&�!��>��>��:6ʸX6D���u!w9�?���̻\�)\�C�s�
�O4��Og?LV<�%N>��N'h�g�߷~��e�v��z���r�����_��δt�j���ѿ��k��{�3|3n�AX�ƽU^�Vv"���3����V�]��s���c<�k
}��KJ����
���mS�Xe<�Sm[v�������1�@�����o��o*y]!�[�}1�������z�t�>37Rc\w9�\������(�a�?s�#�^%���p��NM�`z`�^}��4�7�
Y����E�$�InG/+q���{������ż����}��[D��0��n�k��٩j�̟XYg[QI�P����g�Y���0\�?��a�8 �V��A��tɻ�ʐ�F�'�e�b; ���'���_����� h��������C$�^��B ~��q�j�.bۻ�Ք%⿒'q���b����0=!�:�͈�uÍX�3f
�/cz�������PK��'f
7.�O�I��Ne�{�睄��^��1�K
��[�Ob?���rY�y�f��р�^�cf�S�2�P�K׎�|��� 	@.�)� /,頗rs�H�7nnzÞ_T��x�R�9?C�3����?o.��aQ���s;�m���'�s`n�5��^�;#�Sz�R�M�%0��6����ju��ԩY���䎡�N�8���$�����i�OY�2�י<�ܪ�tr�x�m}"�_���뻛���(��+2�q6�/c�G�,f(,*ޫs٣Xo��V�w��6~N�uKDO�Ɉ�N�Ldy�J�v.��:��g�y2�^xm��=����I+?/8�z�V�7�F̦:\6�+]�z��I�+ngZ!K�y�ؔ����	1���-VIĽ�zgߓ��^�
���;R��0�@�i���1���X��8xDq�s�ڋV��B���D(�#��.�������I�6����	�b���]I�:��ͬ��f�8��{�R�wZ!��œ��.ǅ�����u�й�n�x�Ϸ\����8�� ������ۏl���fy���$�*�#8�)f����9v@"b@*�o�!O�1����O��#5��1o��i"��u��$����ˤ�ݰ��a�dzr����n>���!Z�ި�����M�R3�QV��G]�?4kS_(���M�j�q��ᴅV^����<��
l��jĉR)���!���#���C�8�.��%L������lԛx�-��p�cS��#���.noHT�B�C��U�b�YS��oփ_$�#�.��
�&�'$Y���).��$z��ʷ��T�7o:�*I��
�O�������3y�!��Ε݈��C3���EА�ΦXy�]�Mï6�S�h�Mw�u��Y]g�8<��aU����N��o����V���햑f_S�A�F����&&�|����
ͬ���F�\�b\�H8�����,5/{�{BW�s����6)��qT���:�����єO%5|�Ge�Y��79`�R�!�\A�d�KB��{���b����N�ɠ�=��l5��T���g��ފ�Y�ґ�)��3_"hO��^��mn�����+G��FJy,�������u
���g���s�R{�7L����
�t�0�z{�^�鯺��K_�G��4��}y0�'�D<�ˎ��������'�a�$V�z��t�����؃nr�>��f��RBap�	 �����
���kO��Y%�����
S���e��(g��d����*zM�����bB�oʢ�E�j�+�^��� �_`zov�ci�� �/�~���z��b-2��>�����)p�}���Z��#&������|i�&��}�\�\�y���褪�D�bX�;�h�ܩ��=���*�P=/NU�%�85K�0��S��e��f�H��9D�Lϝ� ����{��'�Z  3;֪#Ѭ�����`Q"���/g���w��3cL/�����_r�<~��R\�e�0�ݘi��i$�f���hj�+`ˏ�s�e���_o�V�c����M艪0]z����Kۺ����O�u�xa,Bk`��N4������eYG9)r�����O=]�@O�6LBgD�e[~�JTR��E��6�Z?b3��ωˤ[Q6�h���O�t�4���]Ė�@Y#���!Q�&9�I  �%�jaz��6k��#��҉�E�j���O�zc�g��݆ j�Z�T��Y��������>��n(�53�q�R�yn��:(����E�U�U����hmo+��#S#��G���4�X�fG��	�ӛ09sͺ|���]@�������|��ܯ|�/�!E��Ϊ8��돕�6�h��U����҃��i.\#F=��aC�<�M�Z=@��j��⩂�K�/t���i?-W=)���pW�$[P���]��~��[}��Ch�[}׫P��o��`�����'H�ѯ��Y��v��v�A���y�u�nT��eq�ճ��-��.(Cv����$���᛽�5��݋���GG�ۤ��^��HaNd��_�o�?��JfŊs�!�Tej�\,���I��Z�(w��hl�A����B;R3~�����^�v�OA�o�vB���q&�2R���(�R�CJI;����-� 7|�O*ˣ�Ü���Q�_��Ωv��c�����,V�����Չ:4d�҅�#�1{�x�_o:�k̲18=��=�?6wj�\�1���2��N�8V���?�\t�Ȕ{�e&�����ѿ���"L� �!I_p��}���#; *��)���|�G򐲶�j��1��v�76�{�2` Z̓� 3P�b
���gm'I.~Fza�k�ou$B��˩�F$�cq4����<zX��.~ll�?�w����!�i2�l���Q��ϙ�	8�5g'�8�����^>� ���ެ6�E��-ck>��ߌ�@v�e;{Zz��Cl�2���ڽ+Յ��>Ơpw�:CB�o�E��re�n� 7�6T@�njێUd�5U�Fޙ�^����7��)�ts�Y���a2�5��d*�����M�B�j��L�!'{�Y��z���0M���C�t���ŏ��<��������'����Zr�Rފ����~�N�%W~I,cRZ���<vu%�_W7�m)�*x�^`��h����<L�%��$�'%f����q"�7�H���B�;�-|L�����y,��'r,㕩��g���\t�����d��1O�?s!Q�>.��?�ψ��?&ﴝ��5>�%F�bv`c�M�Qlk�yX���b��W.|kD�FGr�#&���ލi��/��6t�;~g�eUԫ^a��$=�@����Q��T������i���s������Z(���M�Ve�h¶Բ 'fi��-{/;χ�����'ª*"�>�ļn Hك�A_��w�䜼tX*Tg��z���z������_�g@n!���?x=A�7�O5��v'J_���>��P�E�Zp���&B}�Dts���k�X�M_��H��'�T�%]�D��W��3s��}�8"d:
E<��������۬\s7�Wsi�yqq�fl_��[>m�A�X�(v�����U��z��1%�VsN$a+&:�� 1�	"�� Xw���[*�[��z�˿�ds�R|��y1�Ŧ�_�Y�� � ��`�����b@~�x5�=�����D����[צ
�w',VE]�ʐ���Iܩ ���&�]#�,_�M�w�1i�9�α�/��r�-&M�*�ܥN�}DN[�pm�(�<6V��fk��~��gq�H��*sd*yi5�����|�lJf�7�>�f"Z�UѸj,����Bf=s ��W�BT��,h�Ӽaj��f���FΖ�w���bt��P'ܔZL��RӞ���N��z>c)m�q�q
��Ʉy�����_����+�1�d{����Bkn|`z��%s��EM�B? 5H��q-�`?K� ȋ�N�O:{���n3y�J�~bj�`�|?���e��4��ň�A1y����ٷ�K��N�b��s��K�$��bI�-p�Nd̙��ne�(c�ص0�.k�ʩ�� }1^&�J�v��saC�8��o;oS&
�4�:\�P�cAG}�O�4k/����d�s`%vq:��u�A����۲�{��C;&Y�S����Q���+=�#Q<����S��`���Vkz`
���N?�$ɉQ�׈O��S��&i[ȑ��~gd�f���%8	!gl� �3��U����jCT��Mc�����ܰ[m %�����m���]�7�tX��y����E���'>yT@i�0�7~��|�A��J8�f�.!���ηm?A1B`l�����@$��a�����gI���㐒��!����� 0R����?�9��v�f�0D�p��%�u�WfO�	ϴ#�����]gG��$�s��zLs�`l�(a�?�u�F�O���O��b�`VY����$n����Ѹ��H+&�ކ�Z���}�_�\�W5'���a=�r��t+|0#�!3Z��6�(��p�ӎ*�yWW�3��b���}���W��4�'�O�6S�"I��;4z���X���={,�/櫚{o�8?�H8��	"��ЅߑIg�r��.�!�A�G38���ܼ_� ��2W�[��c���Tg�Q6����V��m�B뛥W��%�5���t�uO�U�/��k��c���⦬�A$%���Uc�MA�K���,3���ە�B����E.�G�x���3��� ���\Ȫ�}�Ƞ�3�\�r� �y3�d���6��-����Yd�e�sO]�(���hm�{�"��O�e6�2��)�ŔU���h��>@�AWnQ�̟�Fx�zlX����	!@�Gx�!>������0�?m�.&Q ���ܩ�s�pFu�Ỵ1)d6��N�z�Y���}��l��4�Sg���$)jm��<D ��G���i��w�T�R,��p[�nh��`m͐ф32��<���M���EL�u���A��ـ�xk�w���/TDt�u��� �^b�;Öw�kw_v)����\���Mt�^�I���������$zY.���nz.v�f<@-����-;=J	ކ1A��_��5���k*���ZJ�fx�䂅���x���Ȇ��X�bcdd����[�4hڙ����}���<q����ښ�f�uz�����C(e#������&ﰑ�����	��=���#~3�h�E�i��C���
@n���V��o����2�q=o�.4��p���o{��f��]�Y�0�C�,�BqT�u��8����۵���x(E��"����u�mxhH�HMn����<IH��0�������µ������z�3i���QYުDB�[x|"�*���dE7�P����'�;�o��4��%��	 ���*�@��O�E���/�"ŦO�I�m�1�Y���� v��,>�'�[U�j��!F�${��6>���r.���t`ϵ
/}�q_a���B��>�ҿ���?��k�	ć�￭�5���^i���V�B�Ou6{�v�&�m	O���
�+N&2Fm��&p#���7��Y0@",g���M���G,5������/w}�]74V��'N�@��h.ل�� �`�������Џ�
��8�ۉ>լ����9���P򓱔8N�8av27r	�y��-gbol���Ux��Bs�;�$��cu�Rz8O7H񗉿�*��1�G��I�E�$�=�h�(���T���vlm�{`p&��O;z��b���ٓ���dn
���+S�����jO��GH�	]�(>������.�^N���6
{u�hxk�x�td���Xs��kmx�0��Ѯ�p�����|7z�VdD�DdE_$�����l�u+�����Q�_���DD�,���]/�,�Oy5r�-_�T�:!ظ��������\��We�V�s�!�ln�ǐ�~|C����,���ugj�T#�\�ew���̦����ț!5���O{Y�LP��~��I���G�!d�S�k[)�?o��p^�{��/?�>>�q�>QIf:�/[�G�\)��}t��~I�`�~`�n��}z,��)d__ô����F]-��{iU����4���Ά_/2ebz��A7�����9J?M�������*�&dp+�`Ʃ��$�!ܞ�;��;yǻ�Mfb%����_���쁼��Ns����B���샟�~�O8���k�s�)a�'풻~e��	xE��y�;1�����x��Tg�����z�in1�����b�à�==�1��;�/ׇ�?�0F��E��J��K{��y���߸c��&����%�Xn)��o����{*�bA�M��\uVk�S��_�]2�	�o#�Y������)gՐ=��D��?3�ɾ;��!^��uI)�߷-O��"�q�Am��:Ռ2��P!�@�%-���%���˩k�u�`�cm���Ϙ�ϥ�<EY��������_j�}���џ�}{�����i�74��ĥ�$�� ao��������|,�,X�ۡ5��F�M�>@��!9������\�Eʄ��o��C^M�@Y~�p�ȩ�s܀���A{���Xi�4�=�)@�/�KÛH3��������u��y����"ɓ��ճ䒇L۹�/aرр�Cr��RU�U4$�@�Y5�hN<�7�8@I�yL�y���{y�d�'�U1�� I���||�����	�n5$s[�.��#�k��)Bܫ}���#}�z�s�����\�
+��G-V�#i9�&���q���f����04+��P����ZN�3�{"��|���"P6�gq氎���������R�������0�7�޻EN�%�^h�P�'��-w߹%�J1�׽�E�9�S��1(�胇Ya�j����v��B,��	<��䄒S���Jz�\���I%�xUY7���d�3�� A�Ȇ��炞�S��T�a����"�?C�oo=��9�d�ފ�+��SF�Fc�����u�:!�n>��k����@��J��M���m��!�u�/�\3OW�j��j��.1��F���NbzBד64.�7�'��c���l�
�q-+p�Z��K�)�HŸ�<�ɪ?��R����EP���;覞�������T���q��*��N��O\d���|b�0�������u)���^�|�]��^Ip���|^aQ���r�厬�{!y����Oݲ�usф�mO�� gc��r�`����F�j�7FJpj:є�z��֦�ĝ��<�8�l�d�ťr�*��9���vI�P�@�|��!�8E˨{��nq����Ե��27�=�*QVa��y6���t���yH{��B��w�Jyt;,�B�g���u�����w&�fwE���{~Y�.��΁OIR}�襬��P�	[/zG��f՘�R�E|����q��";�}��'��Mɿ:�d�\|�-�~��}��y��:�z۟'��؈{��߭^8p��K�w$�\�/]\����z���3�غ�E�����9�/�̉qNo�GI�R�Y�er�)wA�^̈́��Yڢ��t���8��WY�MY[ٟE�h��1]؂j_�{�-��S U44n�F�\�+͂8 � )�Y;vU�|��*k!��=��F,/�ٓ4����31���s��UT�9�s���2S�!r4�/������zH��I��P��.�w�B:ݯ���Հe�r1��lF�5,b�@�^3-<f�ÿ	��+ЈO���ϭ���V<������^���2"|�f��F�f���������R��)"����"����A�K	���ɽJ�_�U��A�{��L=��IWh}^j���e��D����J�RVIBHDQ'�I�����S�i� �T��Ff+t
 E���}3���f+@,�t]�Ԍ4�{QBC=�o�?8�<D�xV�ĭ�O#����'�y�7�-a�͎���g��~o��aK�Ŋ6QU��i��	�8uc�s68Ӷ�����,z&��z�S
>�ƌqg}[�N�	R�����Z��^��Z"/b�-���y�;3�"�.F;L \_�m!���*����W}�/�]���X~���_�s,���@M��%��+Ͼ����;�g/���?~�<����M�\�2#���I.�x�Y��n��H<}P�I��XD��Z�$4W�b&����1ݷ���u�DG�b���3��!9
h����
(��s�=?�!���%в6��n��l�C�)T���da��ib�kU=�i�E���W�7O��l�`�'��OC=�-�ID��q5c)N�t"�~�|�b1����\m]�K���D���l|p	ʃAa|�h����{��QD2S)4��"B:�~��Ylλ1�.Ą��Q|O�k���JKG��*�i<3|���i��#�mϬ,ۈ�M��W�4�X7�a�m<�{�����}���8��(�1��*�SݞN'W2���y��m�kǋ#��b���~ښB��g��ȴu�u~aUa}H��@�)�W�Hřk��w2�ˀo =�h�oNw��.�UF9L8G��`�j?x������n6���zmHD�h�Y��u�>�5%��_������8��_��\���4�EM���~S��Bw-��wz�2�w�[���[��/2��Ǎؕ��|/�ѿZ����"z��9��U
֏;F"���Y�ԊC��~xm/��kl�4�Ό�S^V�S߯��"�QMU�#CӶN����*��ܰ8V���emkA)6���r��i�#a �9�WlDg���pg�6�|(E,�~b;ߖ-��ӁPb�&��IX���Bi헍�/2��������[ϬSJ�N�4�gvĮ���
�N��d�T�7*����1cŰ�Y�UWwp����5�	�RU��35C���ǟ��'=5afw��Ĳ�����61r���|+g����!_^*���t�4M,���,����n�d�n�Xz�|O�V�ɧ��g��<�/�ҭR��!X?�|�A���#�'� ���Ԟ��z���!=�2�)Ꙋ`����A���RmII�o0���d8�̟����u��[�!VYF#�K1��"���(�i�*l{�&�Z3�q5W.k�yfY�q�3婸	X%M8or�EN�˅[@N8��K���6�AXY]����;Z��X��#�V-c��>����jŬ!��S�cM���&,�1<M+�+L�6��P��5��H/$�B��mU�%g	�!@�L��^�cD+�f>���*��.ݫTb�0��FtWp�;U��� ���1 &�UA^��c�naa��u,���ƻ�e,�T�%�ߙ�,�
���Ž�.+��Z*�������&(����j�q������~��q58�,�>��~��`�� �Շ<[(���.��*p�D��!sD���=�''c%�H?��P�44�z��m%�����d�i���[Iy�*(��ݳ��u�B��G�넪T�	���p�Q�nH�H����d�ڰ'{ǂOŮ��:�4��G����c�Ŋ�Gi���9i��"*Xy{GM��ى��}�gdݝG��o� ��D������10h��J�Ǔ��6��#S�1�Ƴ�1[���kb)���N�{-��
J ���3��{G:��0"��ܦn	�8� �c� �Mx'q/��T���$���ݹ2Ř���M�%$v�`�����N�m$1�l���=��	�h��7��#bv�XBF�wy�5Sѻ0��͝�
I�^��a�k�3��Ay�Eʮp��dC;3��a�&��}��r�˫
�x�c�<���-5�#ļwv�9 �TW_#;�*��`-�S����/^k�ZKk���<�N�� ��qE�D.������\V�o��w�mC��]�B�(���Xx!5�-$�<;����{�M6_u�K�3L����]xT���0B�-0���̩�[n1ؖ�����F{�?��3��fm� �t��
�hY@X�yQ���ĕl���胟�{��B���{���^�Q����OCIKmzbN+��4'/�G��Dn�#��Y���Z���u���M̖��S����CuJ���Pz�2=�����gȃ%��6�h���D�9f�׏��'9�ȑJ������$����A1��0"��>��N�;�����~/�֚9m+
������Υ��Bt?�	IX�3����"�χ~��P�����\���6ԩ��iL�O�g��zC(20g�1���Yu~�G�_F���v�5�L,�y�Y�hނ0-����[�N����鄰�&I��j�Ο[Y@��l2wB`��$�y��3��a�(W��,c+I{5~ʏ��6ｒ�Fi���Y`kcHc^��`�n:� >_���>qd@�@O�8�r���~燐���a����:8��>�)?���9Sfy26�c*��	�
K0����	2ow:V,�Lgs,.�� ���E�+>�oX�)�7���U;���������*h�f`������P�2��Z�h�bg�N�c�V��*����g'n�3��98c��G����oDX�0��CU�7��%}�)T��3�n���F����n���:$g"���6:L�H|��Z��Ť*�7�ǕsM�ܵ��t�
(G$�.�8Se</��6<P���/��jZr��ƛݭ̦n���K�\�Qo�Lm��z����˘�����)�%=�bu�ͯ{��ǼtR(."�C$�o_�KO�6]�,C��q�'��-�Lt��� ����߄��%1����u'qٱ�efO�r������{�T��s���PL�BF�ل�̧�`���QO�	��B��m�|�s�CJ�ذ��L��)���Ŏ�w��O��%�O���ר���I#�5G$b���������A�iy�T���]�}ߠouo~\��8�h�m�>F��1�,���|�v���!�p�k16�b�0_e���ڠl�"cH�O]NpJXL���m���?�U�G�d>X�oW���� <Pp�a~�:s0��Sr���(^�X���[9�9���L۱����[�ns5տs��~sk�;gT%{m���A;��T�,Ѳ�MgK§��"����6�;s�sS�����G�$�!F��v؎��ՊJʔ�1�(g�� 5I����.lbM�G)2+�+y|o�V �po���M��*�\7��۟�H*E�iCj���n��"W�X�m���
�"<Ey�#�	ˮp��OWG�{��� D��/~#%�k��xF#�M�_�k���
n��g5}�r��#�C�o��6�w���1��u�-,����wJxI%!]�+�p�~\v$L��t��ѻ��x c���g�h6(��|�"����E_�Z�s:�	�$��?b2U{�]�?RyŃ���\�P����i�i�F6�4O%����$���돠<51p����\K/V�c�ep�]
6�p�����UE��nl@gD�=�����1k�����*!Pi
��|prȂ�x�:�ɮ���%_j,�_]��>�-��Лf�rv��Xx��w!/����f��RJ\�����R�GcX#{bs1�F���a5	MHd³�"�������qw>t��Mѩ.�%`(��	m(�b��f.�'�o���� �� o���W"1��Jzey��)ht9D�԰�Yg��y�M�����a�-����/PR��D�%�fQ��;����S)	i	i��A�;E	Bi��;~���w֬�2x�9O�g�S������;��0c ��n���1��FU�q����h���{a�l�bE�#�G
Ctŋ��$�=l�7����ח-�D�D�
Pů)/�1'@l��r�����WpG�j�5=�K���8J�3<cX��v�A�E�I"����#�]c��������\��
�I�g�������'۹��z���*U������v�)
+Z�AG��^S>��D���2O�Fb�ý0�(HM7	�0}�\��f�*�8��3R�]SQ)�Y?;��G�s��>k���]�3��,��?.��bPb/w H8�����3<�K�+��>�4����5T>�o�#I�. ��>��ޘ"�f���Q5�Qղ�{T��.��w��ã��r�hQP�9�9�؈#ب#$nv�љ��B<���iJ�9����=
�L|�?�'�O6�ۗ$E�9�֜�oR.π���]�v�f8��8���
L���~%m.}i;h������*\l"��C�O�%o����(:���X�.~��D�_v�&f�j	�ݭ5�V9��Ƚ޻��T�F���������<HP��  �%pe��@��>�*������J>]��Nޢv-uŋNY+���d9S��J�ʢt.a�I�z�����?z!�H�$+e=߶:3(�R;�Op�!\�
���!��{ӳ{�q�%Ih  (��S�����YM��Ƃ�՟�+�|@G������$��έu�l���*�T�jW��4󣣅�HYR�L%�,'-ʚEo��+��ّp
;\����N����:�,�>��L�?#{��I |'J�;����Bu�q}�����L(�i��){��B��5y�W�fc,E�·F��ܗ�����������AU(6�۸��R�\/�$�y���]����9z��oƮ�ez���o��n�`<1�YT?��QE��~5���BN��>�9���� ���1K�x"A�j�#�B���${�6�·υ�1��>ݣ((�n}s��7������i����]e;�
J�}A$b�Z��pIP�B���ߌ�P=�!��<O2�ɮ�4ߠ�;��,�U>�}[�=��,��SK���=;�=�ɋZ��%�����2��;6��#u�6悱��g��*J�,{�{�E=L�!LGN���"x����H�m�t�kڔ�eˌ�G:L��W�`#*f�u&�\�^�Qѯ��\'G���v�[�+r+��>�e���� �
Y�P4!e"u�d��)��A%��⎅�����u�6ww���2F�F;X݄<���H�뵌N�~��=Uv��t�,��b%�w<����ڠ�.�6֬���v�`H>��_Yjx��w��L$K���?�� 1��O��{�{2d�͋��6䬌�Z�$�tˤ�FQ�0�tD,}�?�}���]�����-�Ϻ�3�/�w���
Oo%��Tfd��,}���e���QL�`!�صxWx`qK%{׭ۊ�l��q_���e���L�t�
�)�����D�Q�L�]��S���| hw ���=��j�k�Q��� �|rç��1�c�J����n\��F��R��y璮��@�2Hp�Ůi�!�I)�%q�f;|�/�_~һ��x�!{{� K������O�� 3�8�%lXU�$#�jE=��N,Q�J�b N�ȫt��[F�a�z�q�"-�^O/L[)�8�ǋ�>�w@�i�@(�J&1<+�r�B��HEǮ��-��/x�?�KU�LQ��rS�?N��V�%6j��o{�0Fp}�%z�\�����$zF��ľ�Vܠm�k��������������CU��o\�*ߕ�+H�۸$)*Q�ꯋ��$�����˚9���Ɔ�l�f�6(/��q&[|W8�*������N?�6�4�R D�q��tq����S	���kL��I
ۜGC'�e��JlWa �G����% 4�,�U�:�Y\��I�,�@r@����������@�ٛ�
�չ#{e�Aj��~B�d��|j�Q�k�Ղ6�\Y6kPJ_�P��~yFH�ӹe{�G�2�|���Z���_��qh����%]�w���	�hw��F�z7GHu�I�+h�o!�|i~,I�h\�ȟ��{��l����H��c�ʥn�s�v��<��Iy`W�/��g�&�P������gs=�"��/4
+���|A�ll@�Ԍ�;26�z;3Cx�ꇓ�����#�(K�\L��<���fs�����eq��t��}�c1<?��,`*�&]1 �IC"���7�X��!����WɉO� Lͥ*|L��؂d�{mtZx�G�Jٸ�����wg�A�h��̡�ރr�\QK�
 9W8#�${�z_d����D�����Mw�Ϫ7�A��S��U3h��E��Sca}\�aP�o�E�?���&���J�[��ɜ��1\�D��G�����Owf �PnΒ��*H���S����N;���:u��+����X'i�&�p�}.��آ�i؞���ٝ�vU�A��pA�*6�&�7?���� ���z=����R�e��b�l���%��O���''�u�_�,YU*��v��L��{�Ԭ��j1x3R	%�j�<�K��^�e�e�����uER�Fu�8]�P��^Y���Q��Ax��.`��4x ��/�1�\d.�ߦ�L����.Z7K�w��w����#���+�)���В���G�=���QdܵЪa/Q1��:�O���Xnf��T�j)',0`A�O� ���8y�y��ޘ�q�˼g�˾d��[;Gq��ޗ� ^�>B9�|hM�f�P��k��3tB,Zj��H��h-j�{PP
��h��������e3s����j|�wR�~���pS��ԏ&���3��-�ŭv��� ;���WzQ<9:É���8!XU� �K���CuQ�E2�7��g�&�v�8�6�~�X(�{�FBUӋxX�q
���f�|?Į�yy5���ǙaX��Vx�7�+&@Sd����
���sQ� ��GR_�����	���$�n`Iq
K��Mc�B,$���4�~��:{��mX��2���S&�s�A�۔���
���1TN��d����so
�]�1;��6�	�ڍq�{^J�v���:L��J-7�V�z��/�QП _v)�{��n���ɂkH����Ҁ���aۋޠ?m���#I
��Y�CX
+���f)>n.pk��="� ML{B�8�z��{0\���LϧS����%���S���!g�-rC�yv�(�P���|��m}��p2u� V���ԑk���%��in�[Mb�>~[��:Z�x~�)V[��vO����O�#Ab�!F�rv̷�AɽNe��,�5	3GL\?��#�x����vט K2?H��;���9��׳��Ѱ���k��q�{#w�T�{���w`FQO1yF�����V���A㑕ѓ��� �Mȋ��$��Rx���@r�/�1���]Ɓ�R�/��������O�j�&<,ߥ�th�4Os�ؤ��}vd�o� �Z�u�=����8�X$Z�m�aC��&u&#>;���|a��d��c�
��:XxR`1�A�ۖ�d�`������� �AqX@��\�X���F��5�}�=��2�T�	N_��OtV�&Y�� �C�7�G8?�{+V��k�Yë��.�gp1��o���w�����ʪ;n\�l���>?uD�}s+PS)k�`��d�,x�����s�쉮��ƈ�z4�,o	��1�#���+�d�P�)9�����g�~����!�)O8����
H*jx>0Dc�.������,Z}-����ʐ����o6�3�E�J�]�Bk;8�D��\V��V�xv�Ʉ��oH�f�jI�z�yN�9�@�+��[�:7@�������l�Zꔯ��1��|�*C�#m�v�����IL�P��m��L2!�xyb!�M���L�5�r��G���F����J����֊��G�v���P|x*��<�6F�k[�0��ʳ��"l��I��K.�ݙ9�7+K_|�4"�
��k��o��L�R���%-3��0��]�V-k9m�C
2;Q��/�\~��'���DE��Gf8C��$��٭b{��i��.e{��8�%f�<?���j6��4u�^�n^��c�E���D$R~�ణg�˹NQ���C(���}.�6�4W}����u�'�^r_��%�����É�,�=+ً��n���:�8�2STN+FQ�tbW� |Ұ�g".�zQN�%��>ո��ȧ�9�X��ܮ�Zvq��k&�<�e��0�ɷ��.X��`V�_C�'2��6��]O���@��8�����n��g��U��)ʹ\jg�9�߻SZ-�P����ެ�.+o̅���d���Q���Գ'�#��;���N㲕h�~�gΐ#���ί������b6��D�S��� $h|a�E��O�e���/� a��S��Vh�ِK8��<7�����E{��Y���z'֐S�ū��7��"��졆�v�)�s��K5���/I�1��T'�6��߉k6����0�~��s�V�˹;�%
�🨜t����p���vv�O�xJ���^���c�z����A���w0c4�O�~,,i� G�֥�Gw>>��aY=o#b�Y]�=�@h���ɚ�0s�US#�y���@G
�'*���D����řK"^P�d+f#�m匷	I�oG�꾿37��l&���:
�|��Us�K���?T'	O��>��DH`��M�W:к���'h�'�Ʉ���w4�=tL�9�d=�G�_��x�c	���&28��s��ñ�N�y�t(O�y���E*�Џz`x���-��l>��C�f��`@	h�O���}����:B����ʠ�h OE�z�K�hD���	����U���8wS0&��˺��ʲ&�������*F��p����{�$����L�o���quN+��f��vYd<��q#g�Z�/#:"�ϳ�K��h(��TM#�������+
��S����>�����酷)�b��t�1)N�2,��|����9����?[q���b���O�|k�/{K�51��\���{���h|�sP�g�I�$��ɮ�=�����
{�u}�G@��?v��N��~d��[S��=�q�'�)��K��&��\8 �K�/����w��e/l�o�g���>�����;(�rǈ1�����E�}\��m+��:�E<��;���Bp	����=��V1)R���&����4Q�Ii\g������Ʃ�E�V9 Uo<R1�8����(Q�ظKsY|�z��e)����xk�xy�c���P7d9���H�*͉]%�R��D��QB���ĕA: .mv#;��n�9��6�4�� �<�R��{	~��X�u��Db|��ÛcS���[��B͵�e\@Q�2t�s���g�e&��·�x���'��`C��!�U���T��U���T\ߛ �!���5��2p�*�1ɗ�R��H^x�X�8}|�Ÿ�Ĩ�i0�3�ҟL���/ܓ`�JP?�se�=�{�_X����[��Kq#L����B���[�����Z�F��,#0����	-�j���4f��!��aZ���_�?�{IC�e0́�D���Q�8�>��j ���5�fl�w��0¬?h��#W�+��]` B�ͭ�>��P��'Xq����Fhu���2���H+�R�,j�������h�b(&:�J��$��������N�>��m���_���h���;������<�^c�=�An�H(�ay�b)͐�[�^8�d��om`T�I#���X��~�Mɐa��\���B��p�&�N����s�<�`��U����P)������S��K[Q/��V銏�V�z�>t���_P����_�V;�����ʇU��=ۭD�ki+VyR���a? =�5K���Q�@lN�-A��u[�0[׉�\(�������\
��Q�&^�����؈��� Xv7N�B��@�
A�:��$�����1�R���c�=xtWg��%�r�����^�[��t����ݽ���G�ي�y����d#�ь�"�V!e���
��MM�_�A(�XV���ēȝ� ���U|�J��w~�k=� 9�b���a���6?�R$� ���o��6�q�4ʺ�O�������,�\�e�r�a\��N�ѕA��速�X�̍3�j*}�7�H	z��\[f���������6�-�_c�,�SO~�-Rm���m���e.��l犱;E�&�~��]���w��H⟸�X7�5����4Y�1Bd�&��5P0jp��{AU�Gb܋�]�pr	Pv�I6Z0�5�p���'�#LNcw����P�0F/��W�/K�P�yI\�=���"�qU|!���!~� ������7^[��,Z��[\ �R�/4�!e#�f�H0q���V{��d0�k��m\��;��=Y��KG��]L�|xU���xQ�m�ty"�J���(�� 6f�n�HL��1���Ƀu*i�Kv�(G�cs&����� �q�,,=���/}��(E�L���2���o[y�0�\H}X���N�{ �e|x��X���?,����0$e]\&}_��jf�D7v�N;����?�.�W�G��"z?e�4<+���F;�!ҩ?Pg���\CEY���9r�#��f���Ҍ9wy�R<��O���3\R#��K�R\m�u�l�ʖ[V�y�~�V���017�����+f��c�������I�z[�-.8�N���4�#�b6ӥ��IJia�jbк�$�<4B��ɬ��l<g7x�6s|+��u�1�ڣ榗#�h��9�X�6����
��f�h�Ŋ��Kl^�����a���qoZ�׺]��$9pzò�V�5���#���=A��:*"���`l�z�ǑfǠ�9��$��o�L+r����&�r�"���$��
��\D{�~X�5��-����*�t���EPa��H�<8=ٚ��#�:�R��ܷA��T�hǺ�[����)e�
^�ɔԑ�%!뱴Z���©&���]�M\|@C���?�}�O{�U�̢&
�粅��� <Wp���#�!�����k(G+y��(�s|�):	�(@����q��l"���0����)��ܨ���G)��������=#���;�Nb|� ��i ĵ#�2�0m[�<��I�������y3eu�2=�ԴI�4�c�ΖND�H�F��C؏�w)䞱�Դ}���F\��N.��֤C^���Oʎ��ណ^"���	��
4�~^��q�q�Q�|+D�)��h��s�}����vE��fpl߳���r��`י��CƉ_.��3�m-��d��&��'�N:��&�!�`Q��p;=`�������J'CI�����ٜ�N���*�y���� ���4j����Ԧ1�>�*�=�����6�"(��c'��[����ӢV���Z.�aIL�ס�����0כ�8�f'[�3��?�6	�@Z<{D���+��S�M�>�r+�l0տ����B�M��J��K1e˝����M��EYs���4����&�ʢ&����w��@HЩ��Ίl谮��N���gȚBH�`;����i�n ��m��_6Ǟ��[�!~ŗ>�݇~�cGg��@�_�!L�d�U���v�Sx������=C��sA�UM����p?MNc�T���N�����Y9)�����~�v_��3�I�<<ڄ�S�I���A	��1݋�k{U�[7���� ������Wç����S��`����wt��p rDG�\b�~��2v�
�����J#�C O
ʭ�+��:'�q�Vb&$W���,�NJ�F������ð"gw9�Y�m�7Ɇ9�>
zM�)�V��u���U(S��m2�j�,���DɈk��#ǺA��b@<��%��D��G$Z�HZ�Al#�x�7�R�MxEbgN������x�o/ rR�ۋ.[�Ϧ7^��fN�ˁk�c�ٳ���g�1ዹ�����7&�ݟQ����V9-���+Q@�~1�]׈��-�ѳ�@@�Ro7����r�i�2x�נM�6��$2�b<��{�naH���)[�Mд�P�n-���.��"�YI�z��Ë�#r��f���c�B�B���ͻI��)�f����o34��:���XH�,����1���_���XJz���~'��O��PQ�C䞠u7�ڠ_�)���,o$��[7b��G1�g-�Bvz��R��lc����V�xă�&�%���t�W�䞡����[���"�!^��(]���Ҹ�x\u���M-Ltu��������^�x3�o�����E�|�E�F��M��Eī]L����;�{��Aڧ4�@�."@�\ʬ�=�!Kh����'��TX��Ż�6R�]�#7U�8�;�7~�A\��!8b��A[;A�[
���(�8�[���L�� �
�Н�+�k> s�*�Jfn{v�Wm9�Z�OJ@� �"z����4�w7���»ΩL��4 ��[��~�Z6�n��Ưtŭ;}<����t���
���	���9�W�A.*�����n�)-���b����(,�g� q��͍��ʚ<���m�����N q6�`�z��!���`��>j;��g?��]e`o/�ь �O}NvM����@d9��Ze��F���N��IU�j�|����?�Q[�����*۰�޶-Y-ڙʻAI�G��/!k|��/G�Z�-�ڽl>{D�n@�u�1��L,m7������^vhHu��*��v�v�aE
x��>�q�� �w���9mN�g�O������v<̐|Q��ͧI
K�2��q{?;3��7l�1�{O=���h���\���9v��{k|O�7R��9h*-�#�Sg`���76Ҁ�nT����������V4�O�`( �}���9�:��OXS	��8�b�2��5��`ʌo�(�V�H!h�TS%�����B9����ڞ/�(�+�ؤ؛�q�j����ɫ��536Fh�=���c3��d���7�E�I�c=�����À�=�|D���D'oF>��<)����_`*k�eO=áP�G����R�'x�Lzd|ʵ����qۙ�����0w#
R����lZع��8�T�e��U�8�h5v��T��l��W]���4��BOĽ�}�ǎ����կ�'������Z���F��W�m�I� ��Z]Ɨp$�|��O� :D�%{�{nW'�s�x;�G0�Kk�2X�N�����]U�G%��n��6Mw�������l��~גcשe��W�ƒ%��⢊��,�Z���X^�}�K(jY�J�M΅n�:ѱ	[p�,ք�o~A��R
� *��-�
\N�=N����t{�����"�� TP�^��kv��Il�/�ftw���?D��J����u��ӣ�|%���ۀ���>šTpAc	����dU}i�޸ӭ���r�<m�VU��|e���n���7�IH3]�U᧖�"K�]W,�۫���'?�����9���~)���/x)-�`��$��"M��k-��n [/��w~'� Sd��dϪ�V�y�ㄾ����{���V�����E]ԉD�O@ʁ�awe1�9w+:�G��q�l���\�%E�mi����J� U���8�BC�3�Pi�����\7КLe�[9�"�Ŗ-~}r��5Vy�E)+��f=_qwt�]��G��X@^�f�^�jԜj�X�֒����_Z��[�a�N��;O��j�H����n�Jp���JiL��a��P1p���o ��^Ґd��v���Y
�]�;1�%���f%@�%�u
=YMHD{�C@l�4���;�|R}��!�?f��υr��8v�k�����z�!������"C���g�?������ג��[智���DG'Yc�5j�N��^�2�z�m$O2E_��pH�_�I~a� g���:�(��D;$}>�QǅF#sf���+Z�
k��po~
�"��Ar�˪Q˥A�x��8�\C?����{B)VJ�d��6�ﺊʷ^�͝�%�̭#@�MTw�2��U��~sm,��l�+���O�nk򿃺^�ߊ8�n�D�'��"�y)� ����	���ӆ�;-�u�?�fZ��'�-_y}L*��i�@g;K���{�ܟ�n<�c,(����g�◖����e7����K��W�əyO��u�Ǆ��W+�vC ���љ��I�Ѵ3�1����Kz<e���*ԋ�=k��TŔ���I��l������fg������O����g.�kch���d�`�$��{}��A.Z ��~#L��
n\� <X�Э�|�2����:�-4�F��a�%��vX�u�F�}�:^��7��}e4��
��z˿N7�0����<ھ*!ݻ!��m� 3�M����ƕ������އ<����Ӧ� ���9�	�J-�$a����%�n^��-2̠uB���7�T[<����Η��L�x(O��]I]�y�3l�h�#mW3�К!Fb�ō@�������<��_���h�,�������/Jͩg�V_r����ԭx9���Wԩ�v�>���t-c�ij>!�}�{�a�?�*�f�����Z��'FϞ����b���QS�6wZ�l��%_�箃�H
�h��q"��EEդ[�xŽ��"�qSl9���?@�sd�w���UBC����������-��!�Ka۟�b�^�k�w�2�>�t�l�b���{�nxލI�t-�v��o.��(W�j,��39��u�$:�$x���3��h�9)� �����ͯ����9W��m:G�kg�6��ԺP�<���g��92{}��V�植���D�.���<M�]�޺DEL��--ɟ���h�>&߹�ǎw�p�|���U!�,4��MZ��7+A���BÊ�^]���h��m�M?"l	�0F�%U������>�l��|9h�bԸp������e�h��?����J3�nSP��5�]��(@��x��j���#�hM��<ǽ>�7e�!Ez��Ӛ�;c�1�_�5�7QN�Xu�Z�H� �EE��D���@:�̒��ć͞���5��Y@/Zr�^��n��I�}:-۰O�cϦ}��-��x�=鿻��;_�"�)�,��6#Ϧl_�떍_���螿��)҇�s�=}�^���2G���A$}��>��`�ǖq8�"�¶?��M`�h���8"�%�6�@9�^1�/�4Z���;�k�h��j��_L��w�3�l�bU���V�{�� 2x���8�׮�bߐވJ�������u�G4"��/��U��WBcԶ��7���{�5��/�"H�7�T�ЊXy}�Ie��ڒCC�@�9?�+�c�8�G��Y��q��Y�fv���Q���b^;)�[yY�.��{�fp+���^K��X�u�W%����6��Dѧ�*�G���l���Y.^. {r�ĉ M�b�}��?&:�E�Z�.ܣY}[C����3�1_k-�b?�;�K\�P��n���[�V�A�Vv��ĸ��B4���N&Zu�xd1�ǖaUx�rd��	����o�8ɻ���/2<�a-�py?���Y�5��|Ļ�/?;���Wm�ZVR�!���v����KO���x�Ͱ�Q��q5���p�M�/�����۹ҵ����Ye���Js�z�~��&�L�������39���c5�u�Y���gU�tĘɩi����8��Ct3�G��ϛ��*�<ȉ����<<dJ{�$�@([��9AXǕe�U��c��<�@��%r�ؑG�#q����NI�T֜��|>�Q����q��S6�K��J�S�op��cr� ���o��q1�8�DpI��|�/q��ԏ7ғ�4o��IT�}ۭ%\&��tt����,⪜I��׏m[����I��$B*G ��a|&^ۤ�s�lV���ͦ��Q����Y@A�o/'j��� ��	3�CB	z�?7sl���I'�d[&(۩|wF��G<��`;��:V�9<v�iQY�S{�;���/$��Z�q�m*0��BH�[G�t��0ǖC�ƅ��	-( �~ ��v<S���P\�Ѕ�vP�#ܣ���ϓ�/P/~��%~��Ǒ�KRX˩O����]��B��j��<���y�����x���"���]���x����J$B���#�H���ͪ<�8akd}�4s��M41�%\�Dg
9�.\�H+*b��8���X��H�G4-�6���NJ2n�����]d�k��&f�.�fv�E-�곿[VD��G.���g�L�8��[����n&���]�55�F�ڊDEPB��i-�ʵ��e��L>������p��Y��&����� ���%�hT�)!v��z�*�?���]��(E0�v��~Ѽ�V|Q-3ؙD$��@�,]�ע+ �-�ዿ���w�l��6��ݱ��h�[gf�ҧ��`�����e��4��6c=Ȋ
�LM��.��6���̡+o���qo����g I�I�y��?��A��=���:�o�{î�a���3��|%K�0ǆx:��`�K%+�\�d��M�gŽ��|P���=�<�f��֡p�\�����'�5��z��J�@-Ng�N7�H�����R��-���h�ßR��B���٨�]����B�,,��ˣ@�M}wD��F�:q��sa��a �3 X��->��e�>����39˓����R�;���9����W�}�D��{A�p����������H�i�������n�^(=y���ސ-o�̭Y��Q�{���x���y� F�s����x1�Mr%��%���xM��ʟ<(?% j��գ��I����<X�ΓulPhX-4��t����N�c��
� �
������Óޞ�Z(>yA�]&�*��ɔ<�O.��c>N���$��3��@B��^�k���
*
�>B��-���Ր��:���n�Mcg%T�h�׍��[��v��%LH�n�E�K�ɠX����~�pCM>@P+̯��(��CF;��������Qh��ֽ{7HY����Y��'�2��)d��ш���n�����jc���r��E���Vld�Y��Ie�:�!���a5�z'�o�6�údg��g̫�]&"�>��ì�6(v�%D�0�!�d��Ja�D�p��$�Bg���������.�	��W����U����nq.�XG�V��s���4�:`�s�8�p�k��
9?#t�n�w��P��,�ѭj��>��e��J��#���y��Y=����M.��S���S1yw��H�����)�F�{| �T��R}���?�~c���?�ǲ�/���QV6ki��ؗ0��87���~�[��ҪP�4˦��i"g�.ũi�7����{Yb����+�q�z�~?��2�j"ˋlqT���Vh��S�u��W��+���3����Q5���n�AY�{���1�ո� ?w �3#\!��*����M46)o-1*�F���
X�M��Z���L���u����>3�-�8��Lr����"PW�|�� ����ѝn�$�vS8S�{-I8�2�� �x�_���\����#�2��OOY�1Y0� b|
�H�Z� \y�:�����ttz����yQ�I��	��H(�.�}���D�7���,j:��֊ǆr��O�[��];{eS8�V6$��7A��U2W������6�N$��nŘD�\h���p?��ي��0�?�!}�L�[�����P:�H�x׻;�4�;zD������k;���{|��9q#�MS��3�:���x^�8��� ��%8Ǝ�?�����vk�tB�����k�Kz�K�gx��?FT�5���T�҇�puшJ�p�a���m�5��3I����ш{)���9;�-ܣBA!%��t����ݠ��� Y�g���̕�_z���O?�x	�@��
��}D:ƀ���T�G�FfpVK������J����J�2�_�Q��:�!"4��2�_m��J-�w���<���.z�s�� ���a�A$��a+�D�iy�_%oW�{�UXr���Q{�4�~U�x��&��sz��G���-�H��#��0y2����|��2��多���hʳ�����ޜ(��x�AI@�>��H��Y��|h��9wX@�S�0�'��a@�`z����b1܂E٪Un����1d�$�l�-�o�A�d��o	��<�eHXc� Đ�}��Z�?63��²ţ<і�8�V}&����j4�qy�ﰻ�
i��l!J�����Ft�W��]-�X���x^��aG�F�*֚��e:U��{�t͹�(��+n_R�ܟu��l��AU��������������=͉���
�ϫx3׎���hb)�A�sƨ�Y�'L4P0A&��Z!���23��G���e�lJ\���"	�F���1������"����"��ϙ�8jB�֋ٯ6ؓ!D=�L�.0��U��Ѡ�����D���	�O�mqt��6z�7��K8�/&l�t���_�=ᆅT��"��^P"�z$?��yX0揕�io�S?hj�Nz��4�1����<�B��۹/�1���F�䱺H�����a�n\����P��i���gG��ۈ;�[PmzV���z���Ŏ�ݓu��ݶ���_���"N{�����{Z�}?~��ea�L��ehs1o�qpr����a:v����Ų�o�*���g�qk�ًY=>Kz���y�֤c~\�	�
IQ��nAiΤoS��ҿY3I�Ԝ��п_�����?����`)��j9B^ReǓN�* ȶ�B��5V�(�+��J�Y�e
Bގ$�Ƭ��y ��P�LfT'���-��l�ꍬ�Ύ�7� į���,i��3�dQԄ��n!T�����4�zЋؓ�yX{�����vʒw�?��y��-�cX����"�߀��C�.�z(Dy)$��}����H�2َ�x9�:��D�s�ұ��n�q�=[�k�,_��ˤU$�_۾�Z:�X��*�b�ē�d��пΣ���*���š�(�p�^jC��Me�Oa��di	��R�iT&�+"X5E�*�ߺ�PE�T��#��K/rH� 4�
��ߔ�ԆF�������+l�.f�C��m&5�3�a�*��/f@0�B������v�@E��:����hM<�"��^0K8 k *�>}<�{s�w��\�XMZ�<�c���5|��9&g��ߕ���&�N��2��^p�	'Ц� z���������~��V����4j#+���xw�R��vC�����o�����N׳�&� {|�>�ť��I��ɋ��@W��L�l1U;��(tyQ���2�*a��U��%��D��'(��g��ťF�����/��$~4G�E:��p�����a��e,�-�����<fԄ�|��_m�A^�����w�y����S�?42����a9��_�?=D���d�m�+�ɨ:�L�&��N��<�nQR�D�<>+-[�����E�WT�u��!�@ ��M�+��E����:�O������In��W��}�,,s��)��:#Aۂ+���O�l1��p�T��x�2O����I��Z��69A��%0��̃u�T���zf���M����T�"��9���K�#t������VX��"!y�O/�(���6��XbK�Mm��[��;a�ō��1������{��b�Xp�(v��Ƙt^���0+� O�/��l�[�D����N�y����(&='�G5C���Ց���yݍ��!#�y��"n���$$�fWǐ�i�+�w@��êt��"N�X+��R�ý-��5��4l��{��y6���\����ς�~w����0>��d���ˑ�{���lb�)�!��%�J�����h��B�Nٵ�P���Gem��c��~_���Y�$��E�[��}�݉FybOa`�V?�����Bߘ98��s�5 PZ"�R�qq��nm:�Q�mS�ċ'�vêx&S���Mr�^��da�����,V����%���;��Ͻ����14O� |@�f�M}1�tE�|�,�y�H�*��3��^��/����~�c��'z���4�R�����q�
Cb��� (@���1TNl|b!��� 0�ώ�����	�H�\����hŀ��b`���v*�K#���v��#Z�?�o[1��������'�OU��Y[u��e�Ye��Ѯ	N�7��uo���� �=����|&9��k����J?�Oꨌ&yz�s�S�񁔌?���e�R�e�ĭ0p-�-�Z��p@�����l��N�=xת`�B֔*����և�H_��,�C*���H��]�&�����虣�C��K6��H ����)}F=_��?��7o�
B/U�����F����Ļ/^/h�$����91�%-8��K(�F6����l=�x51�lBTd��'���cx7>$ᅏkq�U�K�v,�]�{C���"��q��tKU������
�=:�p.�]݇�Cj�AJ㠤�W���oTS=ig�[�>�>g
ɧ$$�d�dQT|)虳^�RX��#K��%1�Z������'��k �\����v��>˃t>n����IC
�b�h��"H2�9����)� d�"I�as�҂�����xVpu���x\uv�*���Ы�o&N��//�[�񞾕��%$=��,�u�������G^X�$���zyH4t�����% m-y[�P������	~���Q�������zU������z�>`�D��XiP��������nP�����;����V�������}���|���;s��9g�߹g�
mJ��oK$G�".�ٴ�#�pN�h��p��gOM��is�T]������Ե�$�:�5����w����L�LMg��X@՛y����j;�����Pa�sXx�E��B��mHFDA.�ފ�+� �vM=@a�sI�#���I�򭰛����9����o�b���nF|qS�O�7K�Z�
��S�00�2Z��Z�z �~� E�$��k���Q�Ь\�NO����.�˯�}�>7+$���B�<°4`��$�o ��M��o���,VXSP�DV5�B�%��B���Ò1Br9� 7�o�=X������"p��ױ���!5`�������C���fe�s������A��h^Y?��m������&v�!A�ů��צ}P'Z#EU.�x|桞G�3��-�60��9�vB�p?���+)jd�PW�!�:ݛk��W��uF�h�F@�3N�+O��Y@*|g~7��$�i	s�8���$�I�[��	�Y����k\�����z���ڀJ��	�c_p�L��&/5Pޖqr
�m�h��ŧ~��Xڄ����Є�ݱ����]1t�%��g��'�.Ĳ��ʪ�+�K���}�vm��LQ'9�����GF�G�v�:��T���z���[I�}��Z��~8 �i<�QR�崙��e�dy��#�Su���p�~V��f��Ż,���6� A�Z�pN����~�ArA7>Q =7���FE|��`��qv!n
�#�)4��B�9�����~+��� �7q.�F��3ā�}I4��ؐ*6��5��c��xO�P-0%�:�+��6��<u]�F���FU�QE!<:M)�;z�jn+���y��P���;�FX�Q����[]�l��?�CE����u���`Fޠf^,-Y��0�{�c������e�?N���=%,x0댊��L ���k���r4����?�����xK:���C�p����2I���Y'l��E?�5� ��42὞�l^�Z��]�@�~p5�%�m�'�t���}V��D�b,�E��
*o
��t�mf:��
��YE��W h	;X�Q3���o=�I@����D�U��k�!����;_Ql��H�`R ���i��
���6{Kߩכ�@�*.���������B+���K龾��e�~�CJ��h9��	����FO�ᕜ;�nK=Z�C�-�����mkbxJ��|ؙ�:Hӡ�z�����*��\��e����Oe$?+�l�������o��{�fv;I��u�^UM���?Ӝ]��?��ݕǌ�z��ϯ������$R-E�Z����p�=��e���ls�y�5��;�^�Ρ�ҧ��.N��H�
�zv��=-Dk��`���p�,�%R��+Ĭ�<����|�������V֡������Q������Η�+:��Ou�H����l���dv���M�0bo0��!��т8�yV����J��?��*p�V؏;]�6��,yR=�~�$N*'�;�w���ʜ��\\9��5��cU`c$��d���O)����Z���1L�YcS:���U�Q3���~�ߥܡy���� r�nSqA���m����G�����)r
k��0��+�f�h�fW�PоE���|����:�U�J��ԗ��zEj���z�{gL�?�8;�vO�A�?wy��D��u�Y�i��߽����L��>���NEю^�B0.�Yj��u��ڮbVZ�4��-��=�ר'0i�b(ju"�������+�|�e]w���)��h�ʟuyင���_͉K�Óį���Ӗ���YW�\�nU�l��Pt��(�;$6<,5s隵#L��x;�������s�mG{�ІE ��[�'��*�`I]X}x@�C����x]�E�P6Z�C����E�ù��Z+%�R�{|���y�,�N�^zZ�	1њ�MŢT���E��~sӃ�j�G&���h��c%�[�o�����S.[2���L&{���ky.؋9lx]L�t?"�ƨ;y�h�z'��tC��^�FPR�[7��TϤX���y�5Q���3�����L��0Z幧��p�o�o���}$!啶�*���TT�R��oG�M3b�ԬK�S����thN������ϷĠ(T�H	��}��	}�����8�hCA�q��'П��f�i��Gz����yV��~�6����8�+��FU%�z���ue�H��K�Ҫ���s鰗�����(yv�����C���mW��F���s�脅%�ORFE�,����(�㬆7���maBw��q7����z~���n`P���U�FӒ�y�w{Ϊ���fc����}U����#��pfߒd�^��8�=�ʎ5W��v�[�I��;�	������x�y��2gf�V�ɗ���R�8��Z�/��wb~�7u����5<D�=`8��Dtmz;0RJ|�P��X7qL�P���/�'|/�x����^����	4�rQW:�#��1�ɻjUhz{�!M�M��Y�G��9Ris��ݼ%�L�H����h�ս�ȼ�u��F�q����JaF�'�y����]p~��ǣF't �3*Z�������6�Zz���Uz���*rHy�4�w9��6�_kN'�O��|����lٛ��n�ۏfzXn)��1�O��ɪ��A_%�l.�W��܀��h���FB�Ff=p˙̜^ҪC�6�>έh���1ޓ�1� a��ne��O��R7?��H��5 ���LF�\lI��㵔��J]�;�������F�箆X���7m���2����$_�~�uD��_r� t��Q�i#�"��3	�9Dc���6>��~�����tN���{gkE�p�X���=/��U9����x|֕�<�����xˎR��i��,Wإ�Z/�s�]��C��1ҡ���g.�R ��q����k]�p��i���gX�9<�{���4�q�����ׅ�����lm�89%��@��׋��?Uv����z�
>c'$�Orj���<�*Á+(#Z]�^��l�2U]f�ːi�~��չ◼��`P2�z�!�N��O�l:�L���s��8?�nR8��*ȇ���:u�(E�b��w�R�&Jw��z�/Ah���]o7��l_OR�_ZD�!۰�5v��x)>��\�^���p���~�����e�������핀�Q�y�0@ܔ�_��v0:(��g-(����Ԁ��Lf<�j����M	��5U��֏��4���*��v�W.r+	�߰S;���$�r�sKE} �,�D"��*��Մ�RWY�<�(�"i_�aUBiu8Ed�c`���~g�1�F��Z �y��11��?D<<7������u����ts�|��X�����w�C�f:z e����"���N9`�j`/���ŉ �+'�ԫ�<]��p曜�#��8�m鄜�-o�ݔb��k1�	�tC�v��J�d�����<��D���V�)i럳yc]ڂ`A�9}hS`q2L�<�콎೴�t,�z���7��`<P�ư|]�C���ᒼKZ���R���d^w�^����H�t��7bF��Ğw���]�2IK[��  扝9�]����6[��� �Z�˝�/4���S���}�U��W��H��#4"�ė��͕�T��û�|�з(�$������[�;�GO��#�e
"i�s:���"FJ�"�`}�/�B%����/Bڞ[\u,��љ\����r�<�7"
J�*��.l}UR�rD�� ��س�=�y��,<��`.a�w'�ƅ|����ƅ1��K�_5��PW�A\� �����[h�Ǎ����1���gO�3JX�ɹj�W6$E���>`��[
��Ww�E� ���C�����1�}���v�d|^��T(��.%T��mc��J�����e���i���9� ha��?�7v	z�΀X&�C�-�ɔ�e��ck�k��V>t���5d��3�c���Q	 ��EG�q$ʇW�ӝz���%:���DW@�٭�"`�r:l�ɚaj4$ٖăh�)�j������T�2���Q�w;��_4�~Й��f%�/h�}��@П�e��e����-���hI���Z�T�\m�O�M�����P?z�X��j��(��ԛm�v�݈�"dx�;z�>��Pg����^��r`)�;��︤�9�]i�.U�i�Lϱ�%e�\٘O���Fb5��ךt��r�Sq�~-0���*_�D��۶W��3�Y6��U�,���,�ۚ���I���	��6)y}���Z-I��eh��~�1Fb�������Ҙ��#�s�1�q^u@����CZf��OIo޼$�(�g��cj���8�qr�]Ʊ=8ki��
�Z�A�����v�xC��Esq
\}��$j58��u�����L�>�D�2�?�~R�p�)_�K`_~�73���iă%e$���8u�hE����� E��ǁ�����J(�9Sx�/��E��
&��<��b�#T�f�`�\ٜsz�:��:��=!��`(����(��GLwP�4����:�*#c�ފu`N��HY>!ɤ��B��
��9~t�;�.�k�#�ux�c9�󘮳��>C��-9�S|�.����\�-��/@�E�{J�U�#}�{�����+}Wf��h;@��l��ڴ��xW�8h�߫���|6����ˬ1'l�} �'e"Q_S<g'K��5~�;�z�Șy9̬�{y ���(�:�ǁ��W���]��LK��b��*,�?k�4'��8݆���*d\(_C�C����pނ
V��Я���`D�:���'M��$vo�l�>e��+���bj�V��럺(�!��6)������`e����i�yl��R�ul�Sӎ�V�ԙ�߫�����@���˅pF�TM�Ds�D���q������#�.�L�u��NOmU�s���$���$�i�;R[�3�ㅪ��G{� H�~}��A^7CKc�4��*W�zz�߷W5�:�k�.5���wZix��;gm����`�[g'��E��ED^��|i��Q#p�A�G�_P��[�9����h~��ف(��z_�i}��NOv]B%���2CÏ���G�G�Ǡ-+ ��+��;�s{uZq�2��zh�(�Mh��g �s�̳ET�]�6�����������?�WM�f2O�5�ؗ�sH�L@К"��mK��𰸝����m_���;�ʹ��ל蠌�2�֛�es�h~��חc�� ��ꟹ�a�aO���b�E�+�9��5���ڮ�:���y\'�ޑ��%@�É���j䙎y����Z��~��'m�J[]��ΏF��� Y�P�?���ۏ��+'�8G����܋���M����b	�S��x��o���q9�vk(2�-ϖ�С���GBКf��RCDCXvxO�#;�aEY�O�Kr�}��HpV�o�#k�:�:U�V[pO�m �eס��Ǖƅ�#����J%ZY"`�3(�a�t�`��k�J"A��١l�iw	��X�> �YQ����юO����~�e�:�͔��m�ܧP=�Z�`�)�t�yu@��#�>�vO���^�l�m�$o jY��Ҙ�K��+_�>����*p��>6����i����������~�#8:������1��̀�PU��cA�Ț������X|��V^�E}\mW���)0��(M�G�	�Ղ<0�$>��oR@n�)�W���k6%6�*��~R��)6<����s�ٕ�fl�D}�h�F|�㺰�@�h�zG�}i�1��be$��Ԫr���������+Uud����g	+S\:��И>i����[��jt��צ�\{��Z�T�&r�*rh��7�`�/��?{?/i
���f_c��'P�r�oX����B��GQ�U� E��f(�u���*�D<�p��S%�o�ωB���;!ʕ���1�/9%w{����5��뾻�H�􌴎��n�����G`&��W7��~�������}�`�u5n����F�b6��*�](����&Z�Ԓ�"�|Lw�1��|��x��Ս�v�'�;Q�^U�|�P#����Mw�ToD�� ��Ӕ�v��$Ym%��Y!��+��A����ߙ�A���񉺄�Wƻm��UI_o��}l(T�>�C����uݑ��f>D�ܧ�S�ΪuT�A�u�JH1����B��JR�O���y?�$�����=��G��s.����h/R�%n?�D�{?��)���
k���_����$.�� �Е7Q�s'_�#Y5α� �Ah���g�4�%�Q�����h�ɷ�.�l�=�&����<U��z/J�
��m{�U֌lg�c�GZ�ǅ��_{��;p\[*fc��Q�R��v��u��断��lj����NKK�4�-��o@��NvM�E�(4�\�}�;o��'��LF'˺������a̤Al�TP�t��T�G�����r�ى�m���� sڣu�y��x#;���k��� mb���"][����9��ŢI�W-������Ʀ��	�:w$KƇ���I�8hIik󈱯�Z���,��{�N��G`�pnt�����:��{�<�,h�=�:Z�6��ȱR����=M(|d�8=��} I��I9�H�xpx��s��J4����A~ZJz��8*|����_�La��V�Er��Y��R_n<Ri �I){�>Gy\V���-��^o�*�1��W���ĺ���a	�m_�
���+�I��;�~�N���y�9�?�C�X�f�=�Gn9�z�~��n��`��r��=ae���'�����`{r<��$@Gq mLxe��0����Z��;��ӫ��T�&>����ݦ��˞��*J f��Q[H
e�*6�	���,�5_(�71���"�)�o5(+kb����i��\k�"���w�^�ڽ6��-��������V�v;�N� `6sJ�Y�� ���<Lu)��i:@��+��Q��m��9���Ц�:V��޹�5ݘ�^�oB��ō��b#�<�&E�:9w/Z��"Z�XUk׽:��_�S���͏έ@�sM�L��;�BW���3s�	j|{�Y�{M2�2��� �$���|��d��#؂�C�u�sA#���09��Rbu~sv����Z����_�G �B��ŋ-'�_B�>�+]�niĭB
Iص���k�9�ClV�o�Wk?!�4�Q%���j��fh��G��{����rc'�`��}����O�K]0��=����aP��<����y�7��7gy^�!�� 1y%�\�>-�X�4_��Qȧ��3!�a,��-w�:��k�A���/�	�~�T�vf����3�O��-<W�ʐ��sD���v֮��W�(AI�ɟ�ɐ���"O�L��z�ܫ��&\k^$�?'.��'�Z|�,W�n�S�յ�7�]��4d��Z~��r�@K���|M��~�^�6i���Z��/dA��mź52���?.ԼQê����g�mٌ����qm��2�٧�!���aUǾ_̟@**C����\�$�E�J'c̅~�Kʿ[K���]�pz�d[ۭ�������Y�`B��9Q��bB�˭�Bv���ٶ{n���]�9�qU�2��������AI�7	9吽YGIGl&��W[,KO�~H�o͟K��,aI]�oԂ{f9n�I�|g�vwEVz�7{��B������L��_Zk��p�ڿ}�my뤤c����^��τ�$�Sp|) h��]�d�����Sx[��L��ϬL4 �ҧ������N�9n�p�t#��{��p��XK��W�P59FS�o��6�u�h���19z_2z7m媧��[Z�O>ӛj�/u�|�O<��(V�T�����Z�~d}��q��p�����L����I"�t�8_�U��]�Z���@��Y���]GN�%sl���06��"{3�^߄�j�V���a�Xz�އ5"�Wm��(k�=y��v0������T�-p3 O���v��y�`'�5R�g�BlN:�� w��=6�W."��-FV�){�*XO�����q�D�lbf���3��Z^����>/q�;���\e]s3nsHlM9�΅pٲ��淩b�� c�持����dTA�S�?�Ƽ�Ė���	Ӻvhn˪���!Z�-�n�D%���1��mtU�u�Ih� ��&4��#2-��,�2�u�M��u�c�{㇉��&��6���o0L�_x���i�XC�{�2���/�N��R/	���r~3ࣵ��P�}���d�����W��l��{y5l�\m�j�0m�ن����A��40Ϧ��.��
~23PV'W}&zH��@�mۏ¢�Ӫrw��l%Ԓ&FԘZ�"�.%g����ƴ�*ή�L�L�@�K$�#��x�[����==��'���Yږ���~}�c�U#�X1[DGuazb�r7����r�gy�hÏ�V;�l����u�V"�o�Qs����ci?v�lE����7-t��,�G��nwz�#ߘ	&|;ezm��\Y	�L��&�+;x���j�]�xhw!l�[��D�h��1��j݃49Q��+���e������[�.��$�u�桬��Gu�$坳tQ���Z˕y�~m�b��#�5|�H���kRu�6Z�^?6K?��ݞ�騢�?���^|�md�rp�J�E=����X�C���@"bk��Vѿ�g,K��ژ�Ə|?�R{�`��D$�@v�M<Y��ªm�Krx��ƐC>�1Ӭ?A�Vufe�i<���E����$�Om�Ñ���x�A�r���\Zܦ�W����n>����������ߤ*É�:ն��Ѩ�H��?�Ý�zUm��(��Rt��/t�ĉ�yH����1�X���J���
6PF��]���2���x}T���`��� )��~�z�;����0�>R�l�6�g杜���ln�U�j+n�ir�??f�����@��=j#�{��V,���c3���Z+׷�����:o���H>�ړA��(�Շ�ͳ����!�">����{q&0�Mܭ_��[Ny�o�C���:k\~J��;4���պG�Y��N�[7�tZ����|@w#)m*��r�ݛ���Pp{�h�%-W����D����S��'В+�"�����(�_0���@�X��t����Ρbl����%�w���k�O�-� �"�-�3G�Z��a����~ֽ����"j�:�SA�tr�����+�弎��Ԧ��Q�B�jZ�]�r�)���k�����B{S�6}LnA�Gi�Oxk�����B�]&@8��뷽Z��C�umƥ�?Ң__�� ���Dʌ�9q����g�{yKTj-��\�DVb�G)��Xa-�9顠�]I��)�9�י�;(��V��y����V��5k"�kr��&���M���,{�}�N�_w�/��d�Ns'�l�# 2A��	:���B�DȤ����\KŌż�-�M�h#�yB��(=Dc߉;6��ɰ���Ͽ%N��������"9<$�����^A�Ԥ�k�5/͕F�3�|�7�8]�w�&��ř�[J��y� �-.���p5���i���(�#e�
��X�7���gT��]&ω����/cB��Bf��5�;Y��>��Wm-�]�ב'*:���1FTG�o����3���}"o��g�D��h�kɓJ��׃y0:tW���Q�?abz�4�'S�hxⓔz'��A��<��(��v�ة[`�r�$�����A��U��	<�%�/�F�����ir�J���e�s��Mh�i{^����Z�F�Dдy2jԚ�_i�$��H�c��E|:���QA��Wo'��i�^F�,�O�	�9G�� �����i�O6FE����w����U�c �S�|�*�$q��Z��>��1*�Ѣ+̙�{{ծ��zD�V@xK��I��15T�6z���},�=#�$�y�߻��i�꘴4Me��w��ô-��sO�P�B|�nX>�U�5��t�����P~1I���m�|8w4��x�-c3'�G�ޗ�N�7u���l��mq�#�
'&9�6�S����Ё�O�n�]Q���<��e�2�Äw��ϼ�4"���s�& syH,�T���f0�4�\�_2�bʱR�����J:�k���90X��8�['{p\�Ne�z�����e�L�o���8��<���4�E*G�sV��������(u�)���[�w�lA�-���-��LF�j�	N�B��9�XRcK���f�ފ[�b��?iD+�0�-_���zfA�����UI�c�ެ���^[��X��A]f��@p��Ц���
�4̦���A�)�Xx�6e΂cAT����*5�q	h��T�]��!d���XH1�W�v2�����0Ya9�ɾɃ.�h;4���ҫo���'�h0�:�;��#^\���5)��MۂzV�L�Q(B]'����xD�|�x�1�#������	�F���Y��3z��y\�:��m_��4�APA���9I6��\�IW{�=��(o��.-VM+���R�v\k�9��\�Z��^�� �2�9b9$d+��d\A����X�����ō�o�ac�V�2�`Pr�q�f �0� (�@�z�$p��
�
��Q�2�Œ���k|��O{Ik∬�IcbD`R��|����S�#����n�x�y������$g���K]��J&���6x�[���u�4����T
�����Z�;�w�It�6�� �A��R�F7P��c�o&A|���T����	�����f]�m���L��+<���T��jX�lA�f^��#������f�<6	�8 ����Z`h�j��U�:�lj���UZc���'�p��4j��W�XUO�D�S?�-A�L����=;�L�Eᾛ�0,3��6�5����Z����%D��Řf�Œp'��r�{�7XR��<*�I�C��"h2��Ԃӕ�n��)��U�����y��8$`���ܦll�=�_��ᱏ}�L>��ne�ѻ�	cnƾ�����8��x������� ����p�FWA�nS9�`������%ٝ�LX�G����}5�i8�-|`$���>��[ƾҒ�ե,�	�G��?���WB�f���b*l����:ړ��&�)�����zܐ2���-�2�,-���:��(*N�qu	�\g����B��H�L�F	7���ŗ��9P��&�c*��е3�T��f�	�Y�@�^�:⛄�;��W�b��^E�8��:p�q*:N$�/���)�C�]h���參�S���EL<�-�ŗ$n���k��j=v$%D+�ٻ�S�
��=��N_s��?m{���f�^���[���c�&������O*�b��>ߖ%Ռ$G�tކ�,��Qc����i�T~�0�W�݁(�%�p���B�KX(���yg�3vJg�ތM���U�ݬK��T#,� n���}�������O�ӟ�sw���Sf��C2G �1��
�l�G$�FS+��O��E��N�^i<ݨ>kF��M��Xp�.�K��J�b2a�:Csӡn��Qt�-N����e���������(a��ME��:��e0S�K�_J:�u��*�P���ք�N��o���3t�� 5���`���V���9<�y�Hӈ��vwӫ�	2�AD0|9���]�i���+]�a��E�I��B��3s,����
v�i�|�k>��`.��\!����P+�g���(%&�r{�іg-%�xG��/��g���ZLR^"3(�c��-���r@$�^��Mm����� <���
P����)��㎬����3��vN��}�y&�5ϵ�Ӑ��M�E���F8�����}Qc@ �B��2B#�_�p��
�Y����J��B�ѩ/Q�J�b�F�x���W�'��=�������N�;�筺怒wR��v�Io��p��t�:�Lf��N*�Q��8�x!j'��ʨF��ȳ�.O�E�A*1�U޺�N�s���9�K"=�y|q���[_$D\ e� �<����}l��u��N�2R
څ^�}��.K
�͛�v_��b��y˅�O���D�_�QA8�b��)�\�*N]�?����#���Op^4���w/�]>�Djo{��.L�S���p��	Op���O��nlK8���/0o>3؍fOM���Jvק3f�	;^	�!m��W�/�
ڂ,�HY�Y�#j�t_Ըel9D��2����h�kN&�՜L��w�v6?Q	��s�<�ƽs:z�A|� �X����%c�BC�(���* �D�GRc�<��^�����?�w�q&��1M�NH2�nסƽ1,z�O���I<�)�@�^�.��.�琳�4愰���I�v�K��f�!���r"���@_*{<��?�����dH�r{�ɣCB���֐AKf��W��h���/*"K�o�S�3��(H�#��ˀ��P6���vc�@Ғ̕�Ӟx)���>,�@����~�<á�`��l�k{I���D��-�g��`���(�P9�vF6��h�7� ���S�.����rc����O���H���b�C�$���*K[�"�����ǕE�����u Ӊ��ȼᥩch}�$��ږ2�� q�dΏ�udz	��ȥ�f�S{��i�������-��W.��@�n.q�fv���RM�۬���C1�?h���w�	|%& �� ,zd;��i2�ѕM����n�U�R���X>�D��>Fb=Uh�=���T����`�ؗ���� طv��ٮ�4�� ��+��X�|�ˣ1���`t�)Xf6s\���Pü�ʋ�#�)y�𹭋�����gx9%��Q�m�0Tv�D{�/� �f�ʡ�����'��B���z�,W s~�0l��ZdǅO\���k��=���q5�i��<��W-�-�I�j7�h�lL�(+��q���]΄���c��+���X�v�l`Ʌ>�e ng��e���U��
�+�5�?KW��/��nQ�>C0��|�+
�i�t��)���˂��M�s�.�I�l�;��b��Ss�=s�	2ro��ף��.|�M�d�h�Bˠ�0Sx� ;��d�k��6a2���X4�2����j�Ҵ���7��q�E�%FJy���Y+�����Sx�N&��Z�{	�b��p@���6k7����E�f0r�/��
s*�<t��:���e��I�ƿ�SR.d�������/E����Ñ� +Ư�/	/�|�S�B�F��k�6�Z��6����d{Lx����`aZ��F��4����֪ܘc�7���E�Ap�D
?.ﲙT�z���J$�`���R�˼t�J�`l<�?1z�����q�Nh�F^ ��ߎ��
�� ���qbR�u�;�K�6������4;��Pᯥ��F�x�����w�����Bi�#�;u.��"yO�y�{e��Q]�O�h�C������r&�}w-�m�	�i�\��-��Gu�i����*7ỡ��u�JS�ܮ�{ZJ���~�'�)/0����P�?�Je@x�����4��l9���Z�֥А"�9��'s�����Sn�I^�[>��^҃�eq���_t�4<C��*�����PD�L�Bu�]r%_+���{Z<��	V�>�5�!�,d���M�b�A:�b#����췫�K��*�X�O�;����iƧ�����JX�{�-`��e�]�_��Q@�0����4~��D	c)q8[�P�*�u!������S��TW���g�F|�-��@���o�t� ��T������N��X
���↥2D}s�
��)s�>\
���̾��C=�\|}��%�S�Q^XB��p �<�Y��1\��*�n,؎N���X�/V�衣͉��{��,{���4I�����\)���38���]�ei���|��%��nr�2x��H𵕵Z��A{
O�)�����ˀ�w�*�VO��Wg����&�S��NɃv"��������Z�̘�H��.��WfSc��#����)F��5�B�%f�Ā�t��V�]���}��3�
�I|��k������v^��2���xh�ŧ�Y�1�M��p�wP#	��P&Y5�5�5�����kR��h�7'�T�K���j�L-yQr�?���f%W�`�M]��B�%G��#���BS�L�����"l��v�:��N����@���ˋ�,�1�w�k�X��$p���l������*̨R~_�q�	�Y�/
�9���5Ш�{�#'c�I�v��V�D6�Nρ��6��SF ��4�AM�՞mi��Өo{5��J�#�u�m�4��$կ��7(���&��9%I�w� �������q>,�&&|F��b����Tg�ϕ�L_�i�ئ�p�TT.��Y ���>�,rG9�dm��Ң|�8{�Q�ԩֻ���ѝ`8��] �=!!:<���W�r��3$��{N?� ��I�ˑ�x�5���<���:�d=�N���o5����2�/�|)Ap�Y���l��8��t8^x�%މ�{��Um��1�;Y������^��+���{n���PF4��J�Z�,��p��a��"k	۸^��n�:(��I�**{��e�(��h>�I���AW!G�^�Gy���>�Z/��ǯ�@��ݱ�4@������`�h�gb�$3��������X.�[�m3�x����%�v�PFTG�l�q�<.�ky�=ִ��	�y���;�����;�$�^N#�:Xz}z�?� ��#Xp��f8��M��Y�ڃ���V�x7	��b��Մ�`�|����1����Z�~��1���ݝO+*��0?��N�w�l�"V2�%zC�	jc�E�%�2��O�&�����
S�D������@�JR�$;��(ٌ���]'�|H��L�y� ����b��GF�_产z�TZ��|�9e��d����
�#�3z18�Ӥ�9�H�1��w��B�W6�~�+�3�4/Pz�CLx�w����g�0Zp3sJ���4����}�^����"Bk/l��cy��b8���ƵZ�A���/t�E{���&<��U������tN�������?�s��x��Ig��@C_kwZ���G�� �_gčYʿu�怶>��K��G�-�b���m�W�*����}$��;:4��@��W[��􈚶��t�����\(t�,�Ew�d�m����](��TNDl��:@@t��"vV1M���p�j-)Y9���b��RQ��{d&R��Ü��|�a??6��t�������(��2�~�� �Cc���%8+�W����K�V�Ñ��������������_z:u�n�f�Qɻϣ��TՆMR�+�{}V�������&�J�1��\\�GE�Q[-l5��r�r����!���F�dҖ��Q��.�!���+�D�ǒ�l�F%�����N�-5��B���/�����D��u�Ed���,:�S��VSw8TǍ�g���K��C��V��?��Rx|�S�ILMKe.��\7���^��M���QM�f����+�D���R�2K�_B��'��@�L�7��K��O"4�/O��?1�Р��<��J�eQ��L%�U��ea������x��c�.-cLO�>�'.�o��}�o[T>(%4H����	�l��>&Ȯ����������#���ym��
�i�9�B�P1��bA$��L�|9�����BN��T��l�k�'A����OM��1,���4�B�=���	��k� 3��|�b�ew�Z���6������(� �ю�Z�XB�&-�������2����"P����G���s}4�5�}�� ! �a5V���k�BEE�)�nx�P{v�_n5���I)kb�o����}���o>���'��7D�>��gz_�E�z �6<���}PSK�BF��r=�9|�b��F��p�[Սӆ+�����2A�0���g��K'E�]\������� # ���.�(�E�u��1C(㶘�?�h]x\V����V������V���kb�o~$����]��j�]w���z�����B	-��<;��.���7P������T� �P��
�߅~��#�s�	\���[/
��߸�0�y����kݰ�ǌ����v��LO�m�M���#M�>í��'�	vmm-�Æ�|Kr惟�_�l�� �T0
P����|�=��+�G�����B��~ŵ�Zv�?|�W�W3Kps�K�|F��}�����}�ٚڑ���7����eB��P��k��E2����S����NI�?��J��)�Z>e%���� P�Ɖ� ~t�_����%ar}���]��'*09n�g 4�	P� w�,�'�J�m?^3\%�wrYͰ��N��Z�%�C�[�������N��{�W�CR����i���L��[�Xx\�IҹG+�� !���ܰ�����$8��p.��J.�S55��{����;���?/3~
>�oII!�k�Jp���%��1��������r�iqII-#\yO�A��?�V�������nh�&*�=����-�}2�x�r�D(��y|U�!��V?%p��]ZZ
蹷���n\��T������0"DI�55οނ����������g�%���B�������_bڠKHJ���EQ���u���#ʚ�_wH
��$���?5�|q�2�������D����E	;@L����kA',� �/T�毒���)g��],�A���O�����>��ϧ����(@������/�Lxn��?�:���[~l���[
ܻ� '8'��ę��A$���#ihP![)�K�����u~��B����a��O�\��f��9�7
�e�O����;Π{�����}��Q�d��D� �-K�ޢ�-�E]��%�A��{�,��������^?��˜9s�����<~�e�o�C/"�-���X������4��k�|�/J�B��Ũ,�7��JJ�9��gsU��Ҥf���F3���1��x��JH�_QB���wK	q|���	)2M�?����˝dm��D���'�?f���.��D���Is�������Q�g�h�߿Ԉ���H��n0�����B��kpZv�F�[޳��fB��o���is2��o��$Ւ"A�Ez�Rq����S��fP��_��A��p�v�x��(J����ui츭3�;��Jo	�7AW[����Z�pm�YlR�_���w�w��S.�n�H�N��~<��,q�K�j)�ż��=�z!:,������}����g��#���F�dkc�J��<�8 ��[���0��;�e]���e��eH�Mߺ�yOi��_� ��WGт��y�K�qkySXo
���R{�<�}U=�4]�~�h�Ϋ ���lLM�6�\�$��sϪjP�MZsi���j?��|���j�ũ�ohP������r<&�A{`���=��A��snD�%��܈hOi�H��&1�L�*ߺ+l�)W���ٯF�t9���I{�rĳzB�����A��E&��qn�H�}�w�WA��յ�E���W��_� � �!�e:��3�|���.ӕ�X��{{��]�gn��;5�Ň�G�4<�p�Hk#H�85�@
���Q�;ɮo���2a�y�ږ����w8�L<x7�6� ғʼpE�������]|�̋+����ޘ%���q@�G%�C���=�����xT(C�㾍�VЈ6foV�rn��'���FTu�~���ۻ�F/�H�%���q���P�+M�<�K�=�m�D��7�`��
rc�ɑ���	|����6"�����@A� ���x܂���+B��Ndf�M�e���-0S�&�'�;��y̵}~��ur�|���"*"���Ot:���	��y7VT�ù����䖅�o� d�*D�{��5R��#DBD�"�F����1��ʗ!اU_|_+��R4pl�����������\����@8���kRE4�n��0OCݯ�.񭣾�l�GV�m ��0`re�=p9�|
Bؓ�>��!F�m�2HL
%`��?������E9%/M���t�>򤷂�u��+��:ٗ
 ,$$�s�_�)��5>��ɀ�l2V�^�f"�PY^%b������K��س�*�d4�٢٨�*�8gr҄@8�.�dه\��[�]=���y����u�B�Dz�/�&׾Zͪ��x5lK+P�~��F��4��r��E]*�C���nTT�t�n��|��Y�T��%�,G�-�=�d8>�c �r��NF`
#@.�.C<�o�	�%�ȓ;��R����c�d�=�5��Fk1�VNA�O��9���qz+���F�̢�]�;����vz���(u��fT�X��
�7H��@����H���gtYs��L�>z��i瀉ؾ�-d5"�C��;Kl	�R�R��9+J��5�7����
Z�����{|���.�!��̔���y�x����.�(���Y� �\Wb����Ӂf�s(��(���@9���a1��!�G�$�|�9��R��[�3?��.��AZk_����Y�H�O¼��f��*:*䇔��-�� k�O
�If�'���i��Na�A�L4�{\�'��Y%Qt��@~poE��:��3?)x��I�6y3baw9p�C�=ȇm}�D ��~~~�{$������4�z�$5��Rs{�4�B�ŵ��Q�FϛO��B��'�
ȡ��G�@��	y��7~���-���q4_cF��n����4�`
���f~�F�͞��tBccc`J�{��� ��n����a��,�T�6�I����׵����hs}	�+	����$H�6��.^ay}s�uL��ī�<3���N3���|�Eq�6a�����'���+N�!�"$����^����Cɯ�� -������}�'*��t�h�д��\bb6�i�l�7@k�Joj�J8�b� �:,"���=� =�@-�}��p��ԉKS�J���̉C�IB������&��_Ά�K��+(+�!(*`�{�Z�f$8@�;}H-����4E�բ�I��.Q� Y4E~'�wڔ��J�	�n��	�N��>����>��������<���"`�&���+�����E��`i7��`ۯ`��L�J0b�����F�\WA	�'��aJ����ׇrpv}s��Zy�ng̦�G�Pڡ�6�P�iA�*�A@�P��_���u�>}�)���CUi��g�÷�[���^�^�C�T���s 9�P�-�h_	� ��� T�����޷��u�M�M�W��9@ľed��*i#�@���������J�ͦ��� �:OUS2�ȇ�ݒ�y<�a�s� 0@�|Jr7(��~'�DY9U{�����٭"
|^�K8F05��*���i^f@��oЦ�e��n:u�dy�<�љl��֟��|�Y�m4�4�ޥ��:C1�q�X�L�D5�\��P�`���g�z�T�[W�!@r��FG	���l�g�o��v8�M�P�_����is����6���H~H�9�. �"�3�e?���m:s��@�%h��.������,H�Y-h@�ǔ��.���X�y ć}��&b� JW��K.�A�nτ�)��)v^ȗ��\k8 D�Ѿ�k�5��K���9���=�9� ����A5G���U /Q B\�%P1%�z������5����d�$٬Z�=��k��ff ��x��FMB侀� � �~�q8ؠ?���ܾoѵ��.��dފ��,�MP��QQ�5s��	oLMeKG�� �������h,���X�:�j��x��V����Ԑ��Y,����V[X��*
eN�l`��͜�t���j�ٿ����>]j���Gx�l�䴼�d��f@��҆���,�i�'� CM}�.W�/�>����5QͺWP���/F� ����U��#�4��U?5���Ŏ�<�'��1� �k�ϼ�<X����.�)l噉��"�2�[ו/ȫ�H>8�(l@�q���Q���AS�Y)�g#������*���T�G��Aw�&S�ǧi�������?��K'�e���]����;�c��e��e=`��v+œK����12߾_n)�L0�_�XI�J�>9T�l4���_pfI�|�jW�Q��-1$�v��QF��Ҵ8�b�tax��[�5�i�P�{�����8|�AɧJt������$����ԡ�K#seIzvm�Ư�x��>�@����}M(/�)��O1¶1]�ޜ����o7�H�'&�''�o��O%�({�,y�Xo���&�U��ﾟ�9�bF����7�W���My�U8U	���؂D�m&�h2�F>D�U�(
&vB���w��*��w����3Z#hhz��3$<�������
�����I�Z374)��S/���.n��\�+�Β&������\�0ooZ��{���w��O�STs���s%��e���>/���ލ�6���Т�"�<}��1���0�?�E ��9A��������T'a���(9k���<K�w	��1d\�;Y�sVY]����M]��l�D�� �\�X���P6��4�Η SA�W� �'wu�;��R���%3��`"RS�P��x��&�c���kg�ɪ���������>~i�������&���͹��M��G��)���6\A�·�\�b[_O� A��+V�,ZT��4���,��ź)UP�{��A����ː��_���i� ��tڼ+����Գ�՞Ʌ�E��p�a�ʧ,���	-|~����)-@�(M9��Ⱦ����;�U�e��`����\�T��ڸ[��I��(����Tˠ����gOU{�~Os*�������+���C�  eQ�3H�_eZ���P.�f�%����H���x-U_-�L��V���c��C�h��7I�S�;g�1�p�2���[&������!�}���_(�/0��a;���65���G1|iP�����w��mc
��]�&'1Ge�#��{�l �M)Tﯶ����c	W@{��MB���Mn�c�&����!��U,M~��fH������ե���eie�lW/�� ֙�*��t��;)���4�c�N ���=l[?w����:zTo�����.�K�l"��vo�;
��.��;�6]�2Ǟ�����B��֒�-G^�%��D� �����l9|!h��u����g��E:'5m&%�|/�ݙ߭�1�Y�D�q�?�K^��g�<n��ta;�S/L%=sg��2�~�.m��hr����N�R���p�l�6L�C!PQ�i/�K�o�:N�
~�u���*|YCPC6�����;�\� �n�{
i�4>q�i�l�e���D8�����/I:�L����$�Mx]�>����s1Z��d�) �����XO�B�32g��oe��:�D�fV�փ���]��!�뾓�=W�;�9R/n�|�� �%=k�6� Hr�M�:kI�0����C��T�&�|O�����l
��}F�^�m��
�R?E��?7�CGc��������[ƪ9[�[ZX.�����Y���ꅸ�3��2�C,���#��wU酹�O2���Y��!�#.�J6�rO7h�^�
�e:.BO�$`��$znș�>��ҕ�tO	���V�L� ���B��l�0��Z�3x�q[��lL�d�@�X�;�FWe;**!6��Uٓ���� �}��b��xM9#�b��m��8�% �X+��&^�+�욇����5`�%���3���O 3 :)�C�G�����g�a�nݭ0�&�Ja�kT��rio2�-~�$��^��(x��b<����|����� �qCA�5>�.�nvӦܵ��:���U[��w�����Q���t�A҆E)$Φ�3Whl�yԒ�c���4���S�&��!��Q�����Ä�P��_X��[`FjF��V��%Zf�>;��;�U.��*��Uw�X��[#�3.$ÐE�t�D6��b��*o�Y����Y������`���Oe@���c�<,�,��|��Ə ��dѥ�iX��{�A�]��uyv��]7h���Ow��N �2���#�qo���˻'�(U�4~
SN�;q�i)z:��2�yn��#�Ӻ���|��9�`P���k�?=9a�N�3�ó�g����+�!g�-���p��9d�]n�J��u�C}��@�������z\4)~�P[9G�H�<�a���;�W�>a���n���0ٟ9�q�P*M�B,k�g��6��B��kh�'���@Y���Mn��1��4�^=p�N�Ae�sy<<�J�UT�>��:�;�8_G������{��%��ݠ��B�*�~���bS�E��P X���8j��Y�U��,<�z�cþ�X�d2r�Y�:=� k	Y�F]��H��W�+~4AbI�/����:�`��x#����rXg;қ}"�k⠀Mo�7�S@�K���ݟ�ĵnr�iu��b|p��4ʳ>c�r$9?�t5�]G�e]m��VH=!���c��%O�h�	@��É��y֊�����=R]�e9^M�<v���]��\�7#���Pd;|o׬�,F�8��np�=��F41�UY�D�*���j���g��.���
'�hi�4ؤ�M��w�p9G��]9d�4=	����ik�j���R�ހZR�:x��{G�@|�f�8�%�������%�4F�% aj! ݂3u��[S!�l��:Y�iQ�$�b�\yp��}���Y���^�Aj�������!��7`�ń�MtzvF�,p�؆�m�q�mb��Cc:�Lc������k8U���)�����ȟ-���4p�h�ǫ��&~�y,��(,H�b���ʾ�����j�4�' `I�d�ڎL���J9q��3yW���U��Cv~%�U�!(ac��M\{cQ�2}�����2'��z�͸�D�7�Z�C�m��u��]I��ݛ�%mu(�Q�������M�����_ܬ=K��FUgх+�<�_��=:��%^O���$cm/�t;ͬ��V�{��H�P���_4T��{c�\�W"���q���&���^@lG��%7Ny��u�S���`�\4�ͦm�a�ĀJ�m==Ӧ�mo{*v��e (�sj�Ϗ�� SK��C���O�4�U�Zj<��g�~���Tr"^�����F��y�L��2m�XY���jV3�x�q�2Fؔj�W���{*�E��M,n-Cȣy0[�n�,M�h" N��])�t`ʫl�����������B��,j����m���wf���g�ބR��e�=4��?;>Wv�#�au�z+9�͉��,�+��{��!)('r����$"k�{#5��Vcj�����
���<#���o�Ql�=_~#�'L'����'��
7�(��u%r�}�G��<���u��{�7q�٧���H[f#����3��k�̀�oI�Ă��uG��P!�z�Pif�S�W��&�~<3��[�3��] 9!�D��h��$�Q^��nx�4�2<���0ĥ��]H%���?Aܟ�R~h6IF�������͑G]����x'󵒪��#�ٹ��v�}ɓ���ݡT�_�Y�%4�T�w�»�Ԝ엿�&6�ik#�ug�f��Rk9 ��qz+�K(Fڛ�K�%g�}~�n��%�d�_�kP`��B�f�\e�]U4k#)#��B@~��r]l����8i���������G�IР�������,g�'	X7��h_D�yo�U_PP:꧔K� �δ��t�� �J���{=z�#�yw��]{����Xq����Bt��"Mµ
�ewrW��,7������H��@�Z2Ȟ�+K����[��IM�3�?��:r�R5���W�E�R�t�h�˦B�*��h�������v0%��[�\ͧ�3>u�GF�a�jɕSJ�se��� ���K �X�������Ԣ���T��~W���yճg{4k�Uv��^����A�*G�)�XȢ}�Xt倧��Ngz�)���'P�6[>5g^�v#62\�m6�4��s�� 5�<�Ȳ��d� =�f4�<5�~.n]�K�����(UE��w2�>|d�!g�'�Q2�Ta��c_N5��>����l��e9yyҨ�n�`y	F�_K�����!��j;�)������a+�2��m6��(!��xV����y�D�Sb�Ios]:�iu�e��b�}�|1\�A�j��������
ф�U}ΆƳ@��C�`�M�?L�쉈�v\��������h9`�le:���I�(c��]��N�L����L��'k�skV�o�~�K�	R�NI���)��DǊ�i0 �����K��pu�s3<�&�7����7lߘ��-�L���{�s�p���q�^Z� 5���
���uIj�_;�'��ED ��N.f@�h�~��[s �n�[/w\�t4�B�&RzO���uv?��y~����ޯ'�Ȣ�T�&��ﵶ�u�-�ѹI�K��`~�F\�\)=� �Kx�r@5J_S>�c����K�����y�5�N�ﴇ-�7}��d��I(R٨�,���3�g�o�'+-��M:g�9)t�Y�X�f��3�.�S ��B��K-Q��f����)�2#uvz��L�<�[K�#��A��x_g�c�97l��	T� G�=�'ג�Ũ�f`��/iz�kJޗ�5�(�N��vE�Gwǝ�����_�y��=���u�#�8�
P&�xc.��3m���"y�/�����ݻ�Uo���FD�>���D5��n�)�j�z���|���q�[Bغ��y���d�z�wMT���Wɥ�`!k�V��X�Pé�p�����*,Ú�'����v���������36��2�Y�O�r�O���FԎ=��ݒ�z5v��n�^sՔF��VU�W�~��B50izW�G�W����Yy˒Fu�2I����]D^WQ�r���0�(��r�ҁ���kv4����&<�ց���쇿�dC@�<AT����S̘�������w�w�R1-��$Y)'��0�'�&\�?!Y�u2�,w�����M~�R�ǧh7�?���ᣉ���5���Y��zHU��P����6k�� ���� �M���.ӫ�6��(ZR����FH�#�4�Zտ��]>,�C�I�ank�'��y�����V���
%�N( �F�6e��:�agj�a�_���U|�P6�?p����τ#H��o�#������4��)\|��%��%zGq$�R2ո�R�fZ�|���1.��:״��#`C�0�������A/�g��g{v��|'����*�c�6���I$�/>7{u��T*!�����1�����!��n�3!���&+���FE�7pˣ��_ߠ∙�A`��yl�:��^jBQE��#lXR	�������w[k6�4b<��(ݝ�-��!:O՛+u7K?樍�<B��iTz)(���u�ED�X$s�m���4�k��� �s��q(��g�D�O��OAY�_ctl�_๧]���,<��K\������1ۼV���q�r��6�-RS�>�Uw��}A����U�g_��;�^8�X��T���E���B�|�yr��U P�� n�2��)��"�A�W�ۂ�����f'�e�?@�ئ�-�O�~�蚮藼��Ʃ�����깷�Ʈ��L�18e�0w��T%47���'_��3��H�d�0kz��4-Rbic��9!�`x{�=e�Hj�pv�.���R�	�� 9c���/�v���c�|Z;��9��̈"���k��Q坦�^��>%��3SI(��f�l����/�T�Md���/`�I�#�R�i���+`�]�G���3�#v���7�5� �?��LGWp�ǔ� �5�EM�~�d��	 �HkM����C�/@&���o���|L��n�aE��i� �&��H�R9���L9�K�����S�:9PD�*�`x~�p���&���D���!�z���,	���ht:�s���_����޳���=��������9 DfK]�?��r�������� �t�L�Ri���X��zϒm��#�(yج�L]�K^v���l�B��l�r����q�AD귌�]Us��>��atX������L���k�Y��v��5d[�I��OC���,z%_ k#�P������������r�F���S���m��Ϙ�ʜ����μ}*�ͷ�17㔋��Cs�������Yn�fy��Vxk1�.���Gt+�4��\iX
*�{qg��l���^��"�?-��j@nߧ�7�}D{��G8o�#�4>Fy�HNp_�H|׌��|�|b�e�Q}SP6��9��FE�$v5@T��,��}��6�1���\�! �/��p�F�� H7�:���1&�����\r���q$=��Z�Ga]j�m�/8yvP﮷�b#���~Rm`�mņ�{j��[0͊ݚzy��>�!�·n�wf�!.��C��R���N�Wg*2���,����)�\�Ʋ�w,�z����w'N��^��C�s�g�C��>�*`�+��,�tښR�@�M�W�����s`�0G��������YH$��hK�Х��a�kD������0tŖ�f}� �w[m�6ӯФN�����\�v��� R��M?l����"K$|2�`�����Α 3����my�*8S0 ���Α����9���r�d�+F��Y͕TԵ�΍���=i��1��������=W���PV,�#����6H?��o�#��Ҝ,�P��>�y	XXw��e�z�٨�\ّy���:�d�S�ħa5�5�!G�E�����P��k4��eGէ��ΤyA=�S�G�ʗ���>�r?E�S�鞋�sEM�`����K��Bt ��/Q��]��R�O(�z�G�7����`�)
�q2����~A���_/,}�>�u�G�G#X9���G�ڂ��"�����>��v���6��H�wM�h�K��٪�?�[��K���a����^�����s�ء�&�pؼq�H�:�ݖ`�1������G.j[\������z2��&� u#l*L�D{�KL����J|*@�4�g����@�����J"��&d��@�́[�Nov/d���
�|4,�y�m�o$��x�;�0T��q��s�	�Q�1��p,�$���@�*��:+���3�N�x9X�W���V ؝#�6��|d���k�ë��'��R$�<ز�j,Z����Lv�58��P�������\� �F�RCѮ�ÏE��?�o�eYg�8���C7X�����H�I�������B#�~q��g�d�C�K�_.��U%�}��_���NCU��v��հ�N	�E���@�ۣ�Fvx��Oy���4a�Ey+�������3_Ay��s�4w��[�~�u����LZ�����}���箔�ތ3���#-�����0���()�uX�r~h|#m�:)��{��yq��*�O�c�Fc2���4b��2����D2�!�Ǯ�N��'��E����B�p��!�V�M�����&7�lě W���)��*�(,�ST���E[=�_ƟT�l�Tpp��JlZ+�h1k6I� �#^%ҕg�\��zjQ��[?��St?٘vp����R\[Q>�n�|����\�ј�
u ��`*c���ǿ���l�xi<���q����H>�4��ʚ]����c�\�����9��!��3��c����ͪ��i�2�M�0�?���(�1�6H&�CC�fksG/ײ*z�|?��a���}l�����,y��O���t�Ip�}���(!ff9*��(%��3	������E�y� ˫d��8��K���r1݋k���%OZ�UL�i��b��ϖ���t;�ˮ����@��t(���%�{���)<��-����W���'=S_�!j��.�uT��-��i�wr�-�}Rya�N������v��;�6 T��D�V��LU�L��;�N�����Z�1Eړ-;���W��j�
�>OhɄ�}�
M�<y���)��wO��4_�8��ᩝ#�X^��>aT�K�]�Qr��Z@T���F�^klA:J���Y��8=)�J����tD�;]�P������-�F��a2ޝ�����޴Ӝ��ڷ-w��K�)/>� �|���Y�	�����9�W���^�r�6[<8��(uh�c�vJ�F���,b�OB86�^��k���Q����L�.��v.}  縐��z��P�>d����,�����g*K�]qJo�mG�m��)
�Q�����T��ޞ��06>��J>&��R?�%�!���eQ}�?W��Am,Q��\%�z������\�BB�ki�g��3�5�t �����LKr��Zm}�;�Ovs8�\�'�tuM3Ҫ(ח)���	��߭Դ�8[d���C�l}(�дI*�z��3K��ы��vuRucͽ���-�Y��9����\�<���m77m��`�^�B��s�����P��o��i{k���~�*� ��Td����&���rR���b"g��J�gfǲ���(ɬ����*/�]�M�sN*��ԔE�HjWg{:z�L�-G�~�<���?�`;M-����
���2��]e��C��$.��J�M2C	V����T^��5�{�6���*��V���ONԍ���騬;�s���o��w)�FC�x	���	`�m��_��OV���̏,��N)�_�gß�B�vo#�T�x���f���&[O0��~`b��\�D��������}�D�!�{]�z;��nָ@�������p2���A�w�\�k�A����'M�jO�сk�����c.{q�1l�gbfX�q��������+�`JP���������v�"����pM$���S%��ǿ%�=D�F>���'��{�9�9M�n��c��{ƒ&_�)cV����=����e���<@����/��E��N�8�w�RNfv�Z&�wT0��[n�;�DսtF����߈.
.��5�sF��DFN��1�I�i��X��gӌ���Z�b�#y
6�1��L�Gt��7���d�^<�2MaW���]�\��(�N��Ɠ��V���=���A���H�Ԍ�t�
,�\������e'�������0�5�ʣ᥌:���&X�T fZ7˵v�mϡa,��nnnF,Ijڮ�s��	����Y�r82	Q����e��??)T�Vh*,O���l�S-��z0�����"�}ܷr"��j�`<��_U����(���[r���p�5y��:���(L�#\W����˔{h����C�r���`��G����<�C��`��.��J�����oB>�����1=}�(�x	������{c)��'
�����-�b�R��A��S.�co�o�N|o�ǁV�佛D(챚�A�Ň> ��H R٘��_J*��II:lM��ˡ=���d�Pt��su�\g���㻃��ݑJ��߁w*C��{���L��~s�k�����uw�m c��YcXKA����ؠ�v�����v=�����y��^���m�f6�s�L�4ɺ#��E���f3�A���gO�6,o.� �!`�R���,��½	��%e��-��3�����I�FYV訁���������*�W���-���-�e��T����j
^�_����mi>�D�EY8]��ɀy5w6XA��
�>A��]ˉ�w6��ap�RtZЯcY^�4<x�nf����<�{H�5�P�?�_�P*�[�o>�D���C�GG�έ���BѲ��=b�`)r�q�3��#�O�<�w0 ���Ĝħ��]R��;�'�l��i�w�ۭ�$I�'�g-������O	s5nv��W���XC���txk�����~�d���Q��|�k�@�}2���Ϻ�󣂮�Q�^�|�w��,T��K~ɕ�]K2��'ǧ�b�?d���K-eW���/��]ǒ�<��Kˡ�v0c�M��	C�"ߦ��q�d\2>Mzۇ���w�K��F{�M^s�����k6���ηs"�Qm�����U��r�AY����?�\ܙ�Ҽ�~�ۓ_P�ևu�1����|La����	�� �y��7%�qt�3uX���$rQm�i���<yI�p�4� &<����I_��5����?��l�t=<�<�Gb��%
w-������:�=�U}C{`4�_�Բ>�)��hŵ�čb?��P��)�#�*��ħ�5l]w\�[�;�:s[�nxɄ̆�btN}�F���t/����m�E�ɵ��Gݺ҂�_�2�),P^�[?��'�xR%2
-��qg��H
�V7�m0�%O�ƥ`R@�U�9Z�@�}0����`���7�Ò�|�=-5�F���{v�ɭ�̖~k7���hH!�.���!~��&n\ b_Kq�ZK/BYB���L��8��+Q(?�GĜ ���cDt䋶�P�V�%3�����������+ o��C=~�i�WT��T�1�j�(�y����|s{;.��jW���/�⤜�@���\��!�Y�<y��G����OO�d�j�a\�=5�9��R���`+�.�H<~vC�9%qG�SQ���扨�i,�:w���$������JJ��=jކ�ŬJI�U3׽�i�9U�B��?��4U�k4D�q>�[9�xʞ&*&+r��K���f�ĵ:� R�W��C�
$�Qs{!��6���O�ǘ�%s��L�6L*<3�k�׾�টg�3�߇/�L�3��a8{+
��qa�O���5�������&�����v�y�#�ؙ$��D�880���"���f�B�\��o�����W�cp�=�e�Z�W]mV_�	���яO������3��T�7q��{�7�'e���j�q�n�Qۥ��Qk~�D�KQ���������>.6-�����9�t	8Ad���>��	>m� mpR�.���D��A��z����CtO��N�Ǥ�O�\Gn3$�.203G�+%2�8vԎ?��X��z�[��iC"-��{��!����8���S^cL�L�A�qk����_�!�k]š�n��.P�C�z���z���bq�؜2C���W��!��"叙͆퇬��g�X~ʨTT��}/m�3����Rd�͢`����g��Mɞ�<���2�4a�%{���CV'*	ܫb�[����#7^M�@���MZB���~��B���3���T�
*9Q��D	�T��+n�����H�����v� yo5L��j�0�/�G���w�ϔ�K5��ϕܵ�t٩^z��fj����>Os=@��`�ͯ��:�6�@�ݎJ��@k7��!=��gփ<^��sKw���J�[í�V�2"	��}9R_<~�V��E������ٽ�ۈ��'���!OK�!�lV�Ŕ<���W�CP)_K��V�]0���lvu/��õ5��H�����_���^��,�ʢ(x��k%qc�G��v(.p~-�b�71�Í�<�g�Diܕgyb$�*}}�qR�RS�w.�����K����sR�֦��pFҠ���wg��̐&�����t�J�ˏ�u��]l���,9���
Z�����;�<3��U���`PK�f���5���S����K��;�ə��*�ǡ�?��
��[f��X ����Q|�Q�oJ7��`����煆,0�'�{�8�R��ge�\ZSx�=f��z�$©e���X�y F�52��RJZ��Ӎ����ږ�f�����L�?���3�X��t�x��\)dI�t=�_gɓ��5�2����������A���_���Jyt�x�/$�h��=���7&��YG�C8�8�Kq�˨������ދݰ�֛ҳ���6�����R�CqaښR�$F�g$&�����q���7���2%[{���Z�;���g 5>�)�k8���l�񍽎�&��u�<|�h�c�j\���yU��7aCm�.aQJ�Ƒ����Gs�x]n]j��Щ����6��ԣ�;G�?,��
'���Z-6kտ�'�\j�z��o��ћ!
USjJ'!��YJɫ��/e~1`���%k^�*:�H|+V_�U��ͻ�د�HB�e�gEz`���Wb�8�%��j�~��� ��f3?�.J�Ȕ��L��L��\�Fd�L��1d����(�?��pK�j��"�\|��"��ֹ��,�m��H���1�@=Q|C����R��؍V�M�|�����t�<��[Ku�[;���4���P$��X����^jv�DN��P�c�� f��"�;�&������g�����l\��#h���o�:ݙ�V�m&���N�L d�A�QK��� ��e��Wjm>r��|!��M��G))Z��4�>�A��͍�i<{��f���&����A����|[��!.�.��A��K��\~�wo��o�[7�>�xu]g�2��~-�ܨi�+۬�i	"��S�~T��k	b�;��?��@ӂ8�j2�`׋j�rs����mtϭ�e���L��ٜ�/�ؐ�2���p.�y��G�OgX�;C@x�X�l��ǚ���&��'�w����"�~_����g�ɒ^'*�v�����d���A[�2��.��b��+�*�t*7�~��>b��`}v��z5��{�|u%Yƫ�G��*{���?-�mu�
����$�{;��ټ&�5G�-�t"��x�Y4\p0��y�ʫq�J�����z�A�<�(Yog`ԣ��B��(��T�Ӳ,�H�|�^�')WA�1")�cA�7��C���d4�tI����Jj�����*a����ǴTWe��L�c�.���o�#7(�\Kg���
���HV�����YC�A��PN��Ą�c�Y��ď���菔{�v�lK�E@Z�5��f���Ή�I>R�d�	 �����3�'�ɻ�ꒇV-P&=ΔGDҔ��N���G�d?-�)�4��?���p"U�z��b1�M6����}�&�}ȜҌ49ى����kwT� h�eou:]��7��� �RE=��Sr�[��@�AR�g$�h	�;�s�}�?����_3�g�?���@�c�3�'R1��^WήW� ��=<5{�����j��wo���g�>Y_X'o�y�ѨN*��1'��(�����q9 � �����,�Ag����'�Ir�%���ξ�ڎ9�W��u{x�G�ue�X�+��|nt-<�ϰ�BE����Q;Vd�eCm~ˋE)y�HG��T�X\`�l��*�鱭�grϻ�+6��\�V8���B?����qr�F�d�|�o���� ��9@��߇�]:���ǛT\���gO^L-x��ro�J, ��q��'�[b7��C�&�"�.��\�S�>�40���@~a���{�Y���Xށ`�X>��R՛LފM�6_.˖����!f����7]������!.�.��;����7���$ٽ��9ɮV�@�	;@�z#h�_9k=H j�E�ع_;�pb�($��b>=�ou`�/H+Lq���s�P��XNS;��=N�]]	ج�g$Tx=�L5ƿU.��y ��pr�V����eʪ��2��_�[�~��3��*���K��Rs G}36������ۮ��h��w�K�����2`& ����-��M�ApEo=�e$��OpZ�����u"����Wj�	������)�w������7a	u�o�@[ ���Lw�y��]�Jf�ChlX�H�/EŊ徜��oS���>(5�?�:f W��^�c\%��R��eX��
��"�[�_�v��� ����>dQ��F_0�o�"���{#��1'�l >w�q��7 ��G}�:ǖ���;�����6��b̎��W*��Yf�՞<9�8�{�%�@t1�ۃed��Y'�8Y���P�䖎�#�,8?�߉�^������>���#���57��T�V�XY�M�	�$������(+ښꗥM~�;���{Ϩ&��_�2�LD���TA�-ࠈ�R��׈
(A���N � �D@��&Bo	$$9o����ֽ_���d	���g�g?��{�~w�ʓ
O�������O�|I �A�3�7r�l�8���i�C����NM�����e�B~9�~7��FkP��A����y�{v�s=��w��%`�Φ@ȑ$��Eo�Kr����� Xӷ�.y�i��r��6�kRN�i�Iy��X�+�e�7������*����i�w�L�R`�����/;���l2.u:3���TedEĢ�D��T��Ϟ��C"�;	qRZ;3��L��/�̳��u\-�mT.G��\© YK�r~��n/hw��7��g��@N`�C�&�8X&kB�ml%-��U���H���D���*P�'�V����R����zO#(]p��[����$�[}y���\K�~^�r|��L�7�{)Un��p|��+=t��餷9� ���P�T���:0�[��ȏ�g$�
�<לF`�����b$�B���ƣK+5*9g@6&à�yl�`�̛��?�&�c�j�R���H"��ȸnN�L��`ou;��n�Ǳ.2:��۩9�{�C��@�[L=�!S�9��tV��#	c�Ҭd�Ծ��,��&�w���-������mo�ٯ��ev�� �$�]�|@�tr�
 N�.Ϭ�g!��/r}�ށ��c��w�ȨG���Q��p$ⱍi���{g���$��Z��c���e�.ۉ����[��*�$�
�M��`��B�&J�Ҏ�h ���3�9�⡿}���$ ��������G�AI�K���W�����
�oa/\���:<3o��l�11�v��
���.C��B���5km����[���=�� ��>���F�����K^}�R�o�� +1�/F��laCkc�y�bRg���8�I(�9���l�Pݚ�rW�:���c��([=Sn�6Lcm��Yi�s�<�i��=�����9��^@'V?=�ŝ6:U��OQ�U.��أ<��?�و��<�����?��;֟�j<��'W�4u�H�d0��<�����5}'.��1��1�{y"�O�,$b��k���|�k��>�Z�t��n���7��}g��� !M�q�(q{U<�s����y��I�������gxRh�Kl�jL� }W�_�-���l��vl�[�Q$W�S^!�m#�	 !���r�Ǡ��g�۵Q��%E��/��ާ��g�*ϨM�I짉:�|����͜,�F�7i�\�џ�7���?N�����l�{�R��8�7MT����
@o�4�dc��f�`w���z���u2��-��z��c��˳̛��̋��~���?�fΟ��%�.����y�鳿~v?C[�ӯ˿K�k�����]!F���]��������ד	:�i�����Ӷr'5�3����<��o�? PvT�n�p�#�[^�+y9W��`��O���3���9�Sc ����r҈m)�d���,�Vg|K'��ũQh#�u�=7�Z�=}�L��\.\�˾�0fh_P�|~���Px��$��4;H�4�c,WWֈo�x��G^�5��WE�I`@�����r���h�d�8�p {ΪU�0��Zm���_$����j(ri�+D�=MAo� ���I�Y�t\8I_�����1�ɳ���JY�;E���x��5��!�����$���X�=ZE�v�3�Kd���-3o��z�H���Z��2t�&���	�C���O����b�����+�l�V0+�� ���\�SF�B�#��5���b��pO�)��[��í�iզ��֋U�ӱ�DS�(�� ���$�ߛZ\�'iq�C��t-Nއ���d�Fr�~t��d('a%�v���L����Y����NūM����Rp��޷ܮ��z,��#
 7N�4Onp��4�9u���х,�� �]/.���gVw�C�%�J}��j�'i;ť5�I#�Uk��/����^ &~�2�#���W�f��K���܀Z����k=C�#��1�R�Ps��U���+ÑJ��ه�ʲB���*��Z�}<U>28T�Hx�#8|��T�����8�����p�N�M+ӄ�|)��� �B���d���"�9!@��xqSZ}��ȩg,��T�?\�7]-�8��}rXU ���������3;��)��&�j����?�<�[��1{s���\�� _J*0sV�I�$˥�|2�K�iM����� r��t����w��Ɯ�@��h�qɮ�&	� �[�g�ɩ*���݇n>X��Lr2��74v{����G�+�^�^��]&�j��O�]��3?Q�-+�����S����-�#��tL�/Ӭe2_�i!G����$���⟾hY̓oc�[堕���ok�����A��,F���}G�����`| u�q��Ә����1��~-Z	��$�^�B�7ǭI�t���:]�ٿ�f�S���K���|��9;�㤣{��r��Hq�� ���/�_pD�z���I#jDR��m���L��4�*������.�CA��~�Bk���/�TL��*�=~�����Ƨ�rt�뿝��83vJ��j�mj�5uR��<R5Lc=m4;lR�������?$!���Ba!#������4���<^bU��}	�\�H[�q;if���t���di� %
V����Y|!��>]���Ÿ�A�m�������?�3ߛ'W��gט��x�J�B�� +�By��0�v�G*�Ւߠ5�e���؟<w�ޙ./у���$�>��;%���B"Ģ�,wnTޮC�J�BH�V��isNUȝ�my4�T<V�F^Q�y�=|/04܊��;-N�����>�ӡ�2����qr�G����۶1�ٴ���&ŝ�h5��\ ؍�hgq��w���|T��r�{���S���g5�ץ~Q:@������2d]��>�e��J�D>��J���s��(��N�Z^}����6����
�-Q
�Z��3�q�L�U@������޻��ή�*���U?�8�bڑ�|�ncy�<ڬW�}	�@�rX�a�*�)o���z���jz/����?MU��^"�,�K,�^[l��k�S���ڧke����ᤷޟ$p�E	eͿ����ᤣ��v��?�fa_���@��K#���Bv;�a�K�Ɗ�f5'��2�i$hc��C������[���5h
��Z�v���_����t�����l����\�E���gل"W��w��Wø� h��%��E�]��������<���|��s���^3; �B+��%dQoot�'��ї@�b����FS�`�y��*f5~�i�.�}R��'�}��vy�_�3@#��Y�킢�^~%�H\i���/�gH��TX<�4�-]!�(u�lUd��Rڸ�w{}�[�k���x�������B!�r���'U�OVm�d�A.�e�-�� �xe���B��e��x�'!��X-_�o�kt��Z�Y�c���u�Z�y`o�`��� �8�
����f1�C8��yɋ�9 ��;ˁ�R�����yb/�aͨ��`TK���*�-M�3��d��I�<�îmvZ�h�����3�����~CYqQo�N��� �qA]=ޢl��.A��.����h溪�k�G�r����s6�m��A���4,E�©'7�/�"�� /2*M��KKF,�a�O�6;jr��M[��z6|?�f���N�{�x���֋���K�~'x�/�l����heQ=�j�\��7��%ɖ���O��ǆ8�?&��Qy�"�ʇlx�y��t�k2��-�IGo��e/VAϥ��?El�/��c_����Z=�m��\�~U/�_qϘV���][q7m���Ў̲8{�k�Pw�wx�&4�8��P��`�Lg�D1�*�
��T�U�Z�潱�7�v2bc+��h��_���~X�tP��6k�]?/����0����riQ�d�$�Ѐ~�x���{�J>��v�������ύ���u�|}Ů���64�w�E���8ei6?��pJ��{����b��PaV}!�m��B���z��6s��k+;��"0�N>.#� 	 ơ���B�wh.��7�"��^v��)��g�gͅK���,H�v:�#��h���D��+���L���6�q�ߺ*��@c��D��k��O��s�wx_҉D��B΄�wӫno��ĚnM}ز~���mX����06]�n�]_r���y�����D�H� �l;�in]�H������[�nܠ��M7�n�;5��{^T���2�ݓ����eڎx���HD��
��̋M�Y����vA��,������͑mQx������O9@@����*b	Ц���"�ʝ�#ޗ�/��ݶ&MƤ�7�����ii�������/ߐJ�� ��S��|���H}�k����G�,���qX��h��7%�JWe���]T��8�IVE�l<�&�T�vyKЌ���M��a(2d��Id��Y�77��v��Q�8��mi��Õ�R��7�.��,�ܝ���W|�'�%�|�y��A�X�6V�x��7�8�sP�K��h�w{8%���n
���� )/�0�O@q=&�:
�-@����$�[��}1N��c`s��U�9:��T:�4ss�jՆ���{G�Ǻ��-��ú!���ms��&|@^z0�V���}(A��Oӆ�Z�9��m�3uWA��f�g&��0��)�{�ƽ��TbE�_a�3�p�_'��re�1��y t�1�_:s����A�"�r�fX����Uo�� jE5o��������e9h�S#�g��=��F����C���t^20�w��a-v�|avư�1�+]X�nZ�X��T��xs�zp��z���y}5bw��̘IGG�eL�$�-|\��s,9��0��M������.���'3��R0�H��T�-��MQI=P�-T+7l&�����[]�}$�	�p
����X<�"�\m�� ^d�C`�	�]��;�>M*�X_Z۬ݸ�#r������'�'~l��^�Ʈ2��Ua�W��6tBK,�ޞ �N_����^�����9'3�ڃ���mJ � @�QVL�K���i���f�{x���u��o�Z��ŽbU��wr�o�31TOҚ\�����W�^M��i�f���!�m��ݧt��Z��o5�G�B�Ӝii�Bm=~�`�"QC�$u���N���lc]�P")��uL�A�TB^���dĳT�)��T�-�ΥB���1k����T�C�)2�;���6H��;��̑�+�<�^r���p��h��h����v���r��E�����-���2� �s���%�4nm��FF^��nh�-i�2�_Bܧ�vn7�t���(��|�Gn
�sȢ_h������w�k.�w(@+o'k�>�@6Rs�k"X"��)%��kZ���P_�#���d��S�7����X��(��<�tT��UYH�87ِ[�Yjs��x�p�	���`4���m:C^L�(�M��&�Y��Q�4VX���2�	zUT�"��d!ğk� 2khc
�3�߸}}<�i��DQp���2�"h#��i%퐛��}�����|�I��$hI����P�mr'��Jb1���1ㅲx�@��*X��%V����o3/� �9hs����xH'�G}��lO�ʒ����������W�St����o�s���,�Ѱ�Qv��es��G���c+	y�a�_��(�"��rO�8<x<|Xz��_J.A2����E�ċe�s��qsxJ�Cs�������-:��NT�{Bi�0x�Q��OF,�؇�C/ �:�ҵ�c]rR�)o���T�#��O��΂��*�*K���9$������q]k9z���������b�E@��M��Ȳ[�z�x��eӉ �	��s���A ��B[h���۝uK���ϟR2d<���F� �~\��^)���z�;Ay��u?Ku�z�!�C? �3�.N��ۿ��a ��t� ������.Izw���|�](l��.-���$���4�de�>yvK��H'�Ұ\N~I� �QN-rW�~���[���C@b������������C���iV߅5������g�H!��� , u�`���0�Pon��k��ɀ���`1lҰY0���6��f2>k.��u1�������퉊��ĩ�aV�<�x�P���?�}�pҦ� ���Y��?v��_���+��3���1��G��G^MXI���T�������"�5<��ƾ]��L�D��M%�훳\�J�i�e+��>ʙ�6�tW��9����M~i/{ۆ�؈B��d$������'-'}�k��99�����*,w��%�}�/��[������@�?%�Jd��gG��#K�Z;<6_�Ϥu�vs�ǁ%�R�b`P��dc�+%d+��G�#r5��M:u^�������p�,�q,��x�+���4yCC>��H[��&MUw3 5HΑjES<_�T�w��}�����B�C�m�G&�c�ٶ�[����װO=����ryW���ۚ�x�O�������A�1�<�`|��8~v��~1��^�-~�����D�C���)f`������p���;���ZX�b{���*�v|�rYHb�w��?$ꈾє���iA[1����~2���J�\߹���u���n�[Ѥ�`o�.��&!>��F�iv�ᙠ�As\�&Ǜ�k��B�������+(]�9����:P�oc����Зh�@�f~=����ģ�%�o��Z��cv�=����K�E��uMJV�P����(a%mO����X�VC�x������v�n�_��)���PǍE�:�:���H��8����`����&U����晉l�{�&
�DS��j���&ݍ�'$�n��8;Al��S<�W�۾�[��Ɨ��2�<�R��*�����z5P\��I
�v��u���Ǆ�ȍ��+�+�Յ���F���*��s/���Ӫ�MW�=���57Rw(���ݎ��X����-%�'p��1��������+�����)o������f��餵�/��,�c�'ʗ��L��(������Q4J�!N-����u����2����\�g?�Rs��4��ln;V^��+���vJb����놯pkX����6�FKw{�
��>t�gmKH��!�K��t؎�ݷ��Ȏ��煛�a��
,���,�
v���9��z�穲�{���
���ۿ^2���F��O�m,+�Z}<��x(�%����N�u�[����Z"˸*�Ãs����,�.�wR����6K!	K�R�������2��x3��?M�EA��rb�Xq���f�q�eL��P���Bw�6���M� xL����qL��T�&��$�%����A�{4�0|�����5t�`��Bӄ�}���MT��n�:
�gꇽ��p�[3��M:OE�Q��&�I$n�4@����aHvw�be5�z���)�B�&?:dhh��x���E�)���N��Yp����L��Z��u	�rTgb�o�j�P ��uf����)����`.r��8%ʿno�֞���Bj���cn��گ?����\�p�ä֝��������WL�9�FV��U�~��+�_F��FF~\w} W��zr�l�Ǳk�v� ��<h�]k���h�I$�z7ul#»� �㎯���	��uV㲫v�]G�w`Z)T�k�sy}���a��+�Ǣ���`t���^��ng��,�}�f�K;/��=>3Z�5���ܑ����2��|��> 6�^d6���nG\Bj���|���b�2a�r�_?�N[b�䴮�/��G�D �a�gޜ��m��4l�����9�{�/7��>%gu�S"�r���q�H H�o�Qc�1��Q9��o�d(S���:�~��d`�Ӷ�ԤC;r�Ј-O���;»rR��ga_
 s[Hji�/�3�}{h;Q�X(�jG(�537�v䗖YϹ�z������Ѣ��e�\{w��ڿv�~���$�3Ia�ζ�����%P	�%({iz/��V0����rc��ά�xmX���"0Tr�pA�_�R��k��_)?��ci�Q�S?��-������rUϊ?QUh�5�Y'Dހ��lYC���kd$���s��r��dM�,. �a���q-���β����©q2w�v�u�b�k�V�L�
vE��a�����f*&@���MJu,�k�zj;յ9�0M�{�,)��\����\�۱q�C�Eѣ�F�ß?�U?`�@�V�VR��+Id��L)��sa������(��NSu�Z�� *�I���y��nL.��i~9!Đ�O�x��Mo5�[�a�ET��w~	/�w*^{�,��m+��v��H2��6��>�'7>2��Wuj�q�����qc�j4�@	<�>��]���v��Q@��ئ�];�YT�/b��X�A�S�Rig�g����`t��
�Uꕜ���Ä��z�ݏ×9W���2�~R���9隭������)rmU���o��l}���rKtg��<�GahG:Gs���e&��,�Rj/r`�~"y���['�M�`���n�pV玁OIh�WH�����������y�O��ʱ��\	�&q���p�ҭѹ��C�4 xP
�O��ј���}(�^�	wϿA��Y��d����6"�sO��So���[��0H���A��K��45�%Z@��e���0�ٴ6kYJ���&fSt�$V_�9�E�K�x͟��RC_,�ƀ��(|J�P�(�a? �m1�-&*����(W ���R<92ݳ�%V,4�_t�U2��T]U:_\�7��~�r떦�!_�~f�'����O�k�d��o����|��Q^����
�7M��@2��1�5Ӂr1�pϙ�X�H�t�ir"�V�AO��&w᲎�)uY����u[A�=�f�{�Q���} />�a7���������aMW��. = ]�ncJ@���_�(���ᶈ��CatYl��em�
�J�N�k��U�� ���o!�l�j��/��;��X5��?"M�ii\�?� �3XwZ����j'��}p���xX�E`9���?k�ܹ�w�&��)X�n��M��i2�ݯi�̝��*ND�#'�� *�v�3�ks���m��ґSn	��/���FC��p�oq1��,����3 t�MF���{}ΊB�zř��&��E&M:�ܖK>�V`C�Hs6S=M�G����K oU�5��z�6����`�"�^��X2�ǵ�ⶴن.�V�%� ,i����E�}�)X�M���rW9>~�-��	���x��2�E#��������J?�N\c�u%y�%82a��c�_��H��3^��b�Ex�� �:\����m��3v_޴��ɽ����yU�	� x|����zz=�-�����S��v4z@���>��D�;�����2б
�_*:���=��̝�����+�ò�����鶖i��j�	��_�!*zR����VﲏP�2$q�.�̿7m�=T:� ��|h����;��<�p�o����nr�VC���B�Ez�k{���YB^�V�;<�XI���D
qj��~�ʡ��պ���{���p��̳�3R5�U.DE��%��fS��t��k��|�DmI�P��;�����hIXT�T���>����}h�2�;���&I{!uh�G��Aַ���Yh}K�ԧ�~ ����=I��?"��&�G���d�-�4�R�1���q����x�
+c���`�e�&�?����=�D�ĠG�@��p�1`x!<	Ċ�K�F�d���ԥ��T�\�h���y
�F5�!B�L�3��޴��23
*�uGc�L@`�����`��6[�]���0W�_���=�{��H�t�W0������1ll�;�/_���Ηo�@�q9�fy��������ָ7��Ü�"�S�6��\ې:�мw�w7	�����@;��8�Ckas�[�ݒ����3���3�ϯI��L�)>�
&�O�f�Q�Z�/*�(�����SޗQ<�����h��ҭ�G}
`�aЭ���٘��0���2���Ջ�$+є1It�:;�����S�L�ǽ�	b_�G!5O ��\�~������;"��R�q,����Xϝ�G-����+�W�fi�3k�|N M�E��/.��]ܖ���R���CO��Gf����(9 
F/��
N��V�1s�u��d��#���πӷ{Z<��>buS����{v�pŸ�ۛU�"x���,C(AG���މ�O�O�2�f;j��)�E��L�nͿ}rI����DZ��{!�i�@��H/��c�[�XE�����8M/�� ��%� �Qt���3k��=�|�����sS�_��e�:6�r(�p�4����9jr9�7�m䂱yiQ�����_S�,�������	�
���k���j�˩����q�L�gd�&~�~~g�՞Y�j�B��.�#��>t����M|���
v-����& ������G(`�c�>J��):F[���_0�PZ�*�,���؛�F����l&ᚶh�;��)��g&#���;p挿���٨�_�_F!̈́���h[#����l�㣫�-P;T,[N:>����l����5�?�.��K�>�Y_���]�|1Q��@�t� p��k9l�c^�1��/�T�<l�JI��������&�.������=���>S�%H���lPG%12�P�؈��&��H�@�~$�������3?����S1 �,8n�0�ܲ6IU�Ӊfb9��nz������s�Ua��|�  ����)�yv���ˆ�������%	�d�]{�3�;KA	43�(���VH��^rgT"z��� �~R[���;$�0.�lB��-U�b
� ਥ_6��+�yc��7Ռd�R�h������Z��1�o�>Q���|��[J+D���&d7+��$����+T:/����d����8nB��=Z5P�������������͕�����t��R�� ���Әe�3r�j^�:���k��7AA#K�ڇP<RHZ����B}���D���!����DY����Nt|ż�a�oΠ�]��6���;����
4�0L�
�H؊�A�c`( �^v�,�kU����t�By��Kmv<�R ����: m,�Z�˻���_�!�tC��������TJC�����/Uz��������N�aUwÕE����e��3�-��s� Zg�8�U��6k�z7��\0�uJ�x��i)Qi!�V+�|I3��l[��.����琵��� m�Wd�c
���S�Sj9�Df�۵Q�]Ŗ�pV���Y2d����ZSս�~��uF�o�Wl��z��L Z�?(F݂p��_�^�
蚄<�ƛ~(T$ض�+��"n�7�HVߩnzH�  �����'g��B�K����2��f��܉�A�w�[�=vn��L*���z�_�F��dT�{<��{ ��(衽9?[Ҟ5��-��'Y�Ga��&(��RREx�)s�z��F���R}��x����(a�>��쇿����+XB�'�e� TȘ[�����[��Vu�[��u�Rjc��k:�Ƌ�@�4��+s�+��}��;i�����o�o]����|�ѡ�߁_�|vu�yLJ@����A�k:��m��_J]�gr�ΙP��F}5<hsCi�D��>�
M��a@-0 �#���zE~� M�1��E����sA�V#��B �'��i�m���-�R��֫�o���꺅�6��s��ap�R�\s�Ԯ^�� ��m�4��l,�"bB2��K�=G��ۥU�fe�E�-P��}ډ���۩GhR[� �0���O\� zE�y3ɠ[��O�E??���۲�%��=��y�-I˲�,�j�4���s�+�<�&���HBT�lS���s�/������œ?Ν�P9+��ab��ZVZWJG�-�AVZ�蝥�{}��r�V\�f~�������{���ƌ�� 07#�f�RzuRRJ�ZzP�F�hM�y�2,{�0�H)�\@(p#f:�n;���k�Z9=�Yڋ��� ���e��G�~L���!
�ا_��wӺ��,PJ�P��G����,�v�^�[���ރy��?���BrZ�2��
�Z�֟�P��l���mH@LD�͗���e�mo��C!�3[�N��/�4���8Jr��QbuW��5G�j5�"kCf����k�pS��cd�(fR��?�<{�gh���e���N�h!�T	�EH/�wj�o\��������ݒs���\�&�a&kR�� Ϙ��I��97�id~tA�CEwGC�Nb�@��V�l�$kp� v�"���RfE�,G�ы[�%�m���l1�]�PI����[�p��85@B�Z��t���ʰ|e��
�����|�DXZ�u#�m3,Ҁ�~)��ï8{�"w>5�����R���M�Q�9$�xz?5{9?	"�%;�~�&��h�Z Vpe�b��᲻ڍj�7瘴����e��\3ɳE�@y���w,BԒ�R�x���n~4I蚥�>��+��T/`:���V��z^,��|Xf�i�� $_�z�6kϓss|����?���j}F��A����nX6h�PP�W-L̀L�n��c!n6w��rr9�ң�I�Hc�����h/�W�lf�o���i�U�
uE�{��F�E(zyy��u�l����S+��-����TK���˨�f�`�?ű�H����a��ͣ�F�z'4X��2xm�>�t�_|�8��J\��ؐ���l�ZY]�/U�1�0���
G�"atdf.�����'�c��4��UN������X����{��k�!Gʆ�m��H�OB�"6x�2�i��\��*��d�V��;\Pr�~�v<����g9�9JY�@���\���0�++�#���rJ���:�;x��a�[S:�C���a>_M�Rf�������Jb��z��OF~|U���h��S�����yg¦v��������G���@��}5>��b��n��^]x_��:5�v3�kdT��c��T��4��S'�t/��]�@����(*~��]o�P����CxS�>s�ϻ����oΛ�-�1�g��o<ۧ�0����D>T���j� �E4���~�)#�o�?�U�dkDs��sp�撞�k�P���.��F�o��Z}�Y�-��n�j�dw�9��
�,>�3�������/W�9�]۪��م�X�#׽O/���;b�A[ �$�dt�ϖ����Ú[/�����S�v���S�"�;��ԍ�} �3!s�X�%9[	�f��C8͕6�oz����@zMl��p58e�ɧ�J+_�9��4���A�u�.ܶu��*%� ���<zLJ�o6�q��-w:W2~�~e��<��@��%2��K�k��uBBnR����_�S�'�ya�h�m��G&�Ʈ\
)z�;In�m�f莗��S�.Vn}Jr�y�#��4�/OF�+��(��k>��}�ŕ���i��v�gb�=|B��RS���5�� !�u���H$���?�c�S��0�t������Y��O(،$�N掅�gVnL�lX�`t.�0L��h��)>�l�37�G�՘@�r5 ��*#(�[YTr2K�5�M����:n.k�ȌҲZ��c�N�3��>u��XJ�Ȓ
�y��1����\����D@k��5j���Y�����klVk��k	�I���h�)����ݸ�T���ݟ�m��ңF���j?fO�� ���o�@Zc��r۩X�z�c�����J�[a����J�5��ğ;+��~p�V�k�~;jF�+�x�{Ğ��e'&#s7��*[�Z�4�_�SS��A��|wʘ6���͠��!=�t�y��X�C��x���?��0��v�[��5F{��,Ǆ~�xV���=K���`�:	g7{�JC�~v�­ʸ!%�gv���^u��[�����6,�k��8 �����Ğ���ck,[A��U��)���O�����<��^2F�0�l����%$Ͼ(�!,�8�O���=T^pK�K��s}gH�Z���b��O.�����`�(�D%�:S� i�v��������P���4����n�ۧ��=����4ɛY��j�K���f3��Js�/s$���y�m� N��(��^��zWZ�s'b�Ѵ��:���Ƹ��$�=F��ba����B;+�����A�Yd�e�}Q��K�lö��H�48���	��GJ��cZ��`�EԐ��p���'oα��\�{�(ؔz�N���0 U��R˜��μ�t��b_�#���ラ7��u�澯���髞�u?���<G,�sk�_����ߑ��5�O��̆�76 ��7ڮL�R��k6��+�Yگ��4M��T�o��ܑ����������o;�e��D�f���qS#�k.���dΟ�b�3ڑ�Nۥ�y�_�9t<�������3w�y�P�]>e�D��o\�6 S�M!z��妹����bS�HO`�����E�~s���8����%�w��1w�)�b�����Ɨ�mZ�MySO��8`����y^�����l��`FcL�؏�r�*��1qj�Dݪ���wx.Tv�)��1�(���/-ӛ؉.�h߿4���Fڻ;%����la͸q�){�C��!s��)�л�v��j#�S��V�Υq|=����5���^@�,X����~Å�z���$�8��̯ڲ:���[c]QV�W a@���s��A�?,ݫ/U}{�6��q�o
�e��mG��ʛ�L�]^9��b�	M�{Ol_����H���kr�k*-�ʟz>�K�)���*a���	@�=��JX�]�yUq]c��oЊ[z�\�\Q1+�����S��~��%�x���Tіz��(��os5�A��ɦ��+��,Z���ש+�.��_/�q����m�sA�t�mVGSyM�Ͽ�d��("�wc�`*/S��rc��mY��5O���	��֌���a/��^2n���n�I��!�/H��Ր�Ǧ$I�G����ξ���h|�	�\o��n�&,�Q�h�t�b+���!Ֆ������E����'"�䃩�L�3�oв��㲫H*�� o�w�_��J!�R�[�2�^v�f=���u(���Pa�&'�����H��1Bͷ�˻�ǌ����������Q�Ʋ����a��QH~	�q;�(�l+��Cr��afN����7w��m��>v���3҄���!޻��) *M�&]��05�-?��,;(4k�E� 
wH������:^�p����W�i�з�0+t��"fu��G�cˎ��O*̯�qa5m*�aNcM�g�ȋ��=���w���x&*�L�
D�jkaIb��DȂ��LK�ݸd����5h���ui?���&Ď$�q�$�+o�G	��5GAh]�T/-�U#B|��Z�ڷ�����D�&/o���'\-�#i�`�/��w���uV��[͑��,ƒ�M|��P�������	�gӃ1Ӟ�$ͭ�g��Wλ�Thnu ��Cۈ��TKm���,|�D�ρ2B��ڃL���T�N/ş��ȑ�i�	����B~�;.�1�Ub@�n�j���I�+s��𼂗�<��n�ew5J�R��%�vgE[���=�r�b&D�?��i��4�rbXeI/R�� &5�(��X��q���}}+���Nl��Q��AX��H�H�����t'�Jz�x�T�Ϯ&P7?[c�Y�C�E4���]R��;��,r���:�$�����7�55Cn4��Ph5��?~kۦ~���^
O�"��p�bv�%-�s�|���l��4���ҿ!�z$�8!"��<���,&B�*��4����v
��u0��m���]tmj���zCvtv�ŭ�b�}X����8|��'���-�@3ԉ�$|�r���ڊ�tr}���3��t� _(�+	���Ҫ�(���t:A�����O�9�C�����v6�����C�ܴ��s�rg��a�W��t�g;��-�sV9-��{��v���?�~pҚz��!�&\�=@�[4��@� ����f���U�1ƭA�E����y��)yf�U�_��-�kԟ돣!䴌"b��gx�qّ��O�s8 ,���n��E-�����*Ք���)F�O󣩳��uߋ���z��D�=g�P���X�^�eI��c8��_��Q.��K�{,��`U��I�@���?J��a�s�1����q�oe��������z�e��9�f�K���=Ml��>��T��(I���9�0��֧䱵��7�A��	��U��F��յToS�RCZjQ3߮M�'	�j�ޯ|��γ�[�P�wYU��ٿ��NJ�����cH�ܡ�@��a �D6��_�.���48�\�9�}��	��]�'N�5f���2�����0���r1#VÃ�>ya��I:k�+�)"N��Y���M&*�q�tT��d��v|6��K/�0	�-ʗ.Y��G��ed��b�i(��Rw���Z� �~3N�A�_�r�VX�h����" ���w&eag2*�iE#�L�Q��L8n�N��I�fUL,�ih�2�P�b��jh�y�D�j�a�8��'������h՘������Y7)�@��G�ֿ��Y��V�H��	5���k��$$�7J�J�5�r+G��n��[�"���T���wW4�foڊ	R;�sSv���+ݧ�YW�0�Q�\L�m?�{��ПB��4�����jg�~;���|3��A@I�R{J�4JMe�3��cR����_uN�Ov���f}#A�\m+g�����^Mc��)��7���Y�u�A��"J�9��r
]SW��=�93WpXiVB��
�[�P�Ț�>{��r-�h�����IO�����2�i�k���
񥤋|U�`���Q��U1a�DH����bþвp��3������_G5���a,.j)~]��/$�8�*����᫦
;�F"����؍�R��������t��_� u����|�|��^������;�i��4d���D>d#պ\�����b�;��ڢ�QTT@�j�F@AzSP�^CDJT�H��B	��H��A� �;�.5��!��[B����ޟ�~�3#�{�5�3ך{.l>[���h?9_��(X�/�_u�����ܤ#�h_b@Sd�(]�C��횀���?���N�8��.=*�:d�e\i�Ю�W�,���P-��Q���r�0�H�	O�	�^h��j��]W�:��-Vu��b2���]�Z�#����A�xm�X�J��je��b�'�"on^r������Z���Ff�\��i\U��> ��M�z�����
���0F������ż��mb�P����L^7SK�%w���Y a+R+���[8��3�e�����-d����<�o�Q�M���M�i� `{�=d~9p͑��su�<�5\���H��}�׸�4h���A~g���$�.���Yr�_հ`�r*�pE�N��͍��3��,��6@��#&w�c��~y��ԕ��7ݢ#��JV�өal�w�]CH;Vw��Yv>�xU��U���O����hY���+���(�!X&��갊�rO��Y�ݾ�	�(����+��a=|�W�s�q��ʹ�<E�[���zc<�c�\�`/�Z�J�7�2a����9��d��0I���n�i3�����gcW~X���B�^�_og7��FY��1��r�K�=��?��u��ʾ���E2��Q���u�ƃ�#B"Q~7���MWA\D����R ��������0�<i`9.�5%�/*��*b+��t���l�Bt�)��Ւ.��f��]�xq�ȒՐ&O�^+���a`�z�M=FJ��*���C������J/ghd®S���v�9O�{y��.g�y�˟�J�\k�x&��Ee����0-�.��޶w�s4�ؠ�N����lY�^� �C�wc)�TLz���ݘ�t>oO6�b�A7+ޑ\�KMvCc�gz��y��3d��geհ}ЪAlcn0	g-/�����@�T��u���(��f33�����^�Ǿ�Җ�(L�I��Bk�T���j���]���]?�P��5������V��ќH�<����	���HA����j�W�k�w��Ra,��j1��X�a!+��8S��� ��t���C=	�[�
�,�?�`������ݪuҘ[��a&�׾@�w��`]+H�ʯ��$��_=7�']�Dvp�Lª���D-v=W��/�S�w�8�'��׌����vSĨvu�],��qUa-G��Mj3aL�<�73*�/E'9k�ߑ��dc�����d��NC���Lv���d�}?` �s�neI6\�͔#� �t�L�b�d�ZB[��Yq�Ap��/V�UT��q"�=�������C���m�v��]�_��C�e�&�&LDX��9Mx D�x�Z~X���GzWͭ4P||����F����jg���w{G��Z+��.$�B+]WVs��9|b�Y_�x�'�%�И��8�.}��:X���k����~pŬX�H�5!��HO3�"R7�>��7���6�eg@?��ܻ�P�<��ݘ�X��$�'�p��7����{>6�:�I#�_V�4�Rn9yFk6�\��+�a	B#���Yr�]�ͧ���X��A�TVՌ#۲ղ�JǊn�uX;���3ڟS`��i�����P�	5t�1c�����r�~�Ӝ���������6��Q+���'ɶi1���=(zܼ�����P��.�Us����_`��z�i�T[]�� ��� �2��'�9f��CsM��?�|��b8:#�i$��x�V6��?��LT`������������Ak\� Q��dw���.�q�3.�0?�D<����MDC��tW�\U�aəkou7''3|����qaP��4���1ri�����f
ȯ�+�eQdޞ"*w��#�tdY�%"T����Y(xd6�Ql��9����n^�݊����uۢj��z����, Z����Հ��n3���i_�F�#�qk�ْ����D�����ڵ�����%u�������%�۬]k�3 �.3�Yk���G���r& ?���=ˣ)���������� �+��A�Kyx�!��d�s��aTd�$~���`�Ł���e��s�S���Rb�̹�/ݍ����ܕ׻��z�h�v�&�,�MDQ�w�I?2sK�Ye'��W�TJS�,M!b��9�/�� �ѣ})ͤ=������Hݍ����a�:��:��u��P���!|ߴ;�^�>k�{�t�w3ٗ�wC���=�X?���ou)�����BgM%��v(褺_d��K��ݝ\��I^C�U�U�2�.j�*��Z\r�wJ2��M�x��p#b�5�Az��ϩ$��C=�g<��κ�*�\���)t�}pT�	G�u��Z5�����-=�n�������m9�����O�[� r�bU�p��ݙ��Z���߷Ȩ�d5IJ�2�pa���p�қ��6��mTyC-��ɅE�Z�|�U�������1]S�w��Ͳ�/}�Gv.Iv�E�$��ZA{��I����"��oϞn���'�F��ES7��;{���#�q2!q҇R��	�$�w�s:,~7}�f�}�кT�},�E�m�a�O��J�m`�'�=����]M�}T��{��Βg�ZV�U�#ϩ��m�y��� �6f���@��H�cs\���uJ�Dn`�a��t;;��{�JH^g�\e��!��<�m�iY}�i���n�)Td�Ï�a�ꣻ�:^�)�yZ�:Z�P+g����
�mWS�M�6L.�)qD�#��ov@��)۳o����d��+uO%nL��[,�2�%؍o;�6��1�����c���!0�����*�w�ܚ{h�`7�B�X��-nL�Q����Ma��:i�_d^���Z�]gvѺ[����yd����dEsl�B�*�GƫavD`�ov@0�Th�4��z�
taJ������8hs�ʊ��~No���Jh� i��ܲm���)�(�	����x����~��s	R��ڛ�t饡y˰M�Y�U-0m়v�c\h�H� uZ���G9���:e��md����O ������e�)R+��*���#)o?g��]�E�8ǐ��ԗ�@=v�樈��SQ��t4GJ��=F5���{kU�X��ON`�6����!�8�� v�» �3�ýGY� ����g���K��k��Zc�(�Pi���,v@r�/r-^T�O�=�~�B����yUw�����2�U�0��o��TǕ��~o �y�if��㦄8�V~�kȨwQ�?p�u��?>z��Sd�T^������W %f��s��T ���Zh���H�}��"瓊��- o��3��]J�6�Ռ�dYƈ� �[~~�%X��+��I۷^܂�d��I��p �1�κ�`ٺ���1qţ������p	䄕��_���\�$_���H�D����/ 
��0���Q��B��%m[^<b�x��>e�����M>�/_7��4E'�j�	�9P������G�F��<; ��i!�h��v��~@�v/����s_��'��E�ӍҾ��q�S�f�@k�,�g��o?7_'u;����	�M��A��Lf.�����}�3��	Zq�;��Z�x�4���y-1���]tr�ps7�4t�$�+�F�(�o��픗�h��;[T�N�BS��Q�!S$-V�2ˉ�(Y�v#�8�����Ig2�G;���h�~���CUF�)P3�9Y˽���
�,���S�|zP������>�w���aZ׹s���*ˠ�HU�_�������ם
���~#��b���CW�B�JЩ=i��tϼ�-v���v|.X�I=c��U��u��BK��
�����	˘n������_���	�44u����%"G#4S\_�_�{�������Ť��-�zn#2�m�co�m�W?�Ο���7>��|.vSZR�/mrF�d�ZZ0�f������E���H���Jk5�DE��ș}�u��[w �Yߞ�n��7^>�����)��y�<N�&;�@���i:ް�W^�R��8i��"�ga"ZZ��Ū��+���ί�.�J�9�=�ٽ�t��H���<�������$d
w�ls�嵅+� ��Q�]��m�o��� ��ދK>i>U���T��G��,�,�J��N\��i���,Q�G�_�^1i?)��5�������%�>4'�v]����0��!o��!~�o"ݨ��;�ĩp�-�x�k��ŠZVנ��7����RN�k	�I���h�'�6�N�.ߪ�5�ٺ�Y�g4�Y�Nr_��5<Qq�g�-!<��}�G�?�¥7{K��w�e^�����|�]�UGSc�#������LK�	Et����p��0�"ή ��K0����&�P���X�
Ҕ�[g�`���"�7c5�i�/?���1[;��J���5;�3��dzP[�S�� ��-pF�q�i�$�楨-��%�z�ԷEG���� ����; ��8��,1��gc%jl��,�H?�|��� _��з�II=F|���<�Q�'�9�َg�6w��jd`U$��B8;���r�9������ g��θ��4�qj"je����!��X���dy -WѨ�s�w��*;ȟ�����֩vEw��2��-�'���$$�Yd�R�����lG�/ĝtY���X���2}n��z_������2v9����L���SXhf�d'�ץ�o�F�A���<NQ��W�S��з$��X�I����%/�F� �2L0[�GV�gC��� Y��혓�(|�xQ�R�N�79�1�� �.�mݎQ��&��]���m�#� �Jh�3��uz%��Xl�ZrAQ��IC-Ȁ4J��2�1�b�	^P��܉+�g^�t~�2K�y���&����	�˸�t��]{�y/ˑ��|����O���X��B.�8����<�ӟ��k������g��7����N��� Ք��_R���:�FO\�X����\?�@SR���Q&����Mg�ܝ��R�!x�r˄��FQ#��K��N�J8ڃ��g��r2��k5��_a�U�"�f���N�Ĺ9'���v\��yP�����Do9"=�n�q�|��~FW�L:cZs?�V/��x�ᖠ~h>o�keUq��m��ɹO�=�Y�|�����Z�'sy�}V�V�G�B���Q0 �ԥ�����5)��u�ӏ�7eջ��I0I5���zd0�z �h��`VOߪ:q�T��h�w*��n9k�	��%<Կ�W�035<�j��ԯ��_Á�a߀?��u��T+[�'��:�4h�6�1?�2�������l���Uc/ۿ i�t`p�h�d� �2]���ox�n���k��I�����8R�@��߫������պ�����������:E�����(n_�o��[t�=���_�wp/�@�f�F���@Ӛ械v�O�0�6�-�r�"#'�
�	�͆�����[�)߆�<�������Pʿ�Q\A���O�'e��ב��c��n{=�.l/�@���"���)P������m���n�ͪ������,��E�'x�ӏ^�=~��K^lp_�ﲅ_���W ���jy�6>'�<�u�oS�so��w8���&���3X@~�a����&
�|$�;�����z[�|��7���zdQPRe����v3��$�����V�k��-fQu�wga�-f���|+��'d�'���!R�>�趉�+�Kg|b�Ъ��w
 �
I��_|"��6��\r����"�C�]���u��T9u=&�߀/���+�c[y�7�"U#�C���#fJP�H�Muc��vϘ�ރ�o��ܭ���$�O�4�<	r�$�Qǽ!��7ɿs�<<��*=)��=9��.~$Q�-]�@��bb?M��s�¯��cƚ������d�z\�{u\R�~�0�+��.� �׮ �LƃF53V�`�+����o���wn�F�N���ty���R4�c
�Uު�w��>�m��@��M�w�Y0�N�4/j"I���on@��<N[�]�\�G���E袞��6Yu�;}�ܔD��� �ڨ6y�d�O	�k��Z)mU ��Ҿ-�)w2Y>��P������>�l+�ક�~���/O��֐g}&Pb<�3�Y�����sG&3�B>bn(�Nl��E�)�~��槽���ޓ��Z�b�m/ݱ�'����xb�A~:`�	����{%���@�t�<��Nq�7V:~��G?k/��w���D��e�9f�q�*_ϙ��t��$ �u�r�?�F-A>�w��2,�����%ɚR3gd.^�%�HO����)��j����]'L�x�g&�]Ѝ���'�z�H�-�]Ht\��݌��9�(Ll���Z���&(��z(w�b��q	�I��E�T^�׳LDys�
5�ԅ�Q��
�	!	���#%z��0�_b�'�O|d[; כ,�u��xdj���ʦ��������x���?��!�~�$%����@O�u�2v��U��'.w�sp��)���{���fO���Īo�K)c��F ����7oU�|˛�Mf�$�!W��X�lchi�A���c�t��y���2�|43믔����=�@��Z���`���W���kݳ�a���}�g��u�y�'YNxԾY�AѲ5�^~�k�-i�����?�9��w�v�Ϭ�kO@�: �W��=��̎��]�6��"˙�����G�X,2��"!�1�`�OX�V�?EX�_�N⮩�w�殁	�̬Wg�H��jeV%�E?��<ޓ1昈��(Z��������LA�.�uQ9�����oD�����wc�^���OZ���-A��ͯ5ȅ�iZ�VE���=���6�\).H)���;�h���!��]�7h%5���σ��[,����i��/5����qu{�&��-�mIK�Ce�.n�)�"�{�i��NZ�SD��}Ql��9���o�Ə��v�G��|�W�~��1���rgݿҟ-���U7"ĨJqH����S��5@�v�ه$�9CYCwme�$N�[�O���Y�W�횬[�ԏ�v���=o�����Jc~�m#�]V֕l	�����΋�qqw�:�����2�j�3��2�w�֯t�n��>O���
ʬ�s<���^í�~�	g����Op�~t$��ڮH��	��>�m��Ģ�a"le"d<O���$>
H-�(=�;T�;�ê%g�����zn~�~b]��x|�ֿ��a�����;��gK�:x�#%��Ͽ�0�D��������OS�^�ZFa/P�=�5ng�
�$Ҧ)��4�_j�'	fe���v����6w���4vz���a��4g(�G�#�ϰ��`����\�ҥK�yv���ҝ��}Fz�<������_^L#�l%3f��F
o�<���e�0ۮ?��H��_{��lF3an�2��r\FtʧM!��0 �wyy�Rt�H��
�Q����z��Kw�is���T��i��ӂ�V�Q�?�ˁu�F]oQ"���Q���@v15,Ǩ�p��3<Z�����i~V��8�����;�����x{vq8:l�2���i�`�&������|�յ�o$^�:TB+t��}�"�sa{��J��i��|mm�$]P�(�lC`�3��Z��ϲ6'$��O�o}��7N���DJ�7���:�w����b\l�3�/�P���oس-��W1�xҏ�v9
QͱiݕЬW:���(��x�_c�GY�|�"UK�۟;�����zf=0I5�i�P��/o���z���K�����m��/�����`��k0� ��<hsٔrJSg誤�
��~��A�"i,���ožQAj�e��U^��S�W��I�;*<���㒦���G�Q�؉�_��P��;b�	M�c��Yv/��?�2�-	#"�&$����:c��n��e�값R&����u�����,qy�<Nx%��;P420S~��ಎ�0�AL^X(7��3!������@��9����^n�Wq�����q �*PD+��Bk9'��̮����PgfQ�����I�Zeߵ�<�����5�4��,]V�/ "� �h8'{��|W)��=`f���RY�1��d�E&���� �x訩#���B���܃y����%�X�J�BΖ���t��є/����hPD���4�a�� ���IZ���"��.���S>�
��E^ ��.Q
��p) ?5��*�7l�;���/~����2���c�t=���}q)��|�d�Ġ����tA��(SX�S�Y!
�Z�/�<r8�^&����X�i�������*��1jvg��j���R� 5�S>z��i��>ϖ�.a3aTiE�꥚�)s��[�[���|d�)H�'�`\�΢��k�G���Ш��F��c��W��T���O����'� �	��?j�A�%����ٴ��a30��%	Uu�)*��}�9|%So�&��4ř���?w����$I?.z<s�&W�:Ҳ2��̭Ƃ
�i��H��o�|ň�s�}D�e*� o�����k&�{��n����${�Ʊf�ɝ�|CY�'vi��,	��c��Y�U�7k�8�)�m&�M����O/�B���ޭ�ϕ����F'y�+�T�₊�QU�[����u�d�>e�7V\��
n�ƪL�:�	Ǡ���I��k8]8Q�N��|dO��ި|��y�r�퇩~��ʩ���R�saԍ�[Mk�xC!_� ��L�O��>�4h�`�J֙nߋ�ս��jU�2p��rƉg ��/�6��+_��'���Q���eq �����{�pQ����a<� �;1|�+��'-<�A������ɷ�Ԕ��
$�<N�i�l����H�$5X�e��:��f��~	�9г�-� �޽�P�><c���Z�����8�m��n��2�Z�x�Ŷ����_Q5��u��1���.U�F�,֍����z�r��V>r��9h㓧i������_
_�u��݌0Yo����ڙ^b����(�WqT﭂_\ �_��_c���jy��Ƴ8�w*��C}.���?���J*�t�S�r��䡋7��ڊ��7>>d�QxJ�
�Qx�isUX6?}����Kmؚ>�>�q	��"��T��nR�
x�y[�����s�o��,�t���k�lu�����Ĉ�h�P�N������ϗjR������&!2cB��W�T��"�^�{��,Ĉ�>5	n;��I�!r�F�?`�\ �w��0�J66w����(W ��R*	�*��@�֓J fڥB���O�Z�U{�3p1s���έ�V8�H��
��l���U=���sn�A�N�g�d=������#��}� ����屋��X6h�>�3*Ϙ��8B}��j��FY#P"��QkX�����d!@��u�ƚ�q$0�,Dw�C`=�g�%ʪ�Y����`cE�4R��� ?�t�r[rH/��:�Ra�D�pW�^j.���Z�:��⥃#�l7H�~˨�D�N���!#������= �޸�'s_��~hq����(�,P��|%rK�D�R�(�mY�N�munq��ߗ3cF�h^��#~�5�^��ҳ����<���t�ƚ�e� �jR�]�M�QS����o���w�]���M�������Ĳ�D�O�e{��]#m�4��T��� ��z}���?ǅ��$	>����w�Aֈ� 2��RIS���U�>AXܒu�]	j�&�@)�&��j��h��h���`n��^���� Ǚ��Z�-e[���v(x������%xX	(`��1��=Q���`ފ�sL>z�q��S�T���h�A����H�e԰D��I��7b����뒕�?��]}�Ik��wӻ����ӧ�����ӷ/��-|PZ�Rx�~����X�[;����ߺF�y�ǭ�+E'dR�W��;r�����xख��U�^���y��M�jj��~��d�kiQѰ�q���g������ ��'�ç[�՛�	خ�G�X�nL�e]�`%]�[~i-g���r/��yy�ʣr0����\�ѺR��f�՗���_<��uh�{36�_�#��0�l�y�ֈ���wo����T8&%W&Y�k�!Y�sg!�l�q�؜�wȬ￝�6�Y������83L~�V���%��,ܛ�BN���Z�ͺ�.��7������f-��PDV���;O!gL?��hZd�]4�O�Ǽ�ݍyÅG�~C�����d�Z�ݠO�f�w�v2��>�lv�p�T:#��$ɱ�Z�%^��?�>|��ȼ_L<!�$���3~[�	�������|�F�1f�L�CXTb��M=_r@�Ty4��������
JV��H>%Y�ty7zq����KLt�sp�2A`\Q_|0�N#�408>*��a���U�T��$�{r*�?w��O���[�ױ�!��ҁf���m�I�������|JWzy x�߉�E�Y��&"
w�x��}b&V�_Th�I��^�:R��Y(�?��M>��*�(�Z��^�X���\���'��&�y5�֕�� |Q�`C.3-���~���"��"F�~0zN8zYHx�y�k36&i��$��}�R�Ѐl.������������mt��Αf�F�X����qZL�V�9�~S�(�'Y��w!�C����k��fק�2ļG!����(�t��ɟg�'j^�`t}}���V���s��I�?�x�뇷�7�����W�1+Π����G�� ��/�f����М����ׯP���HEoi"�?1�I|#�w��cN�J|��j��"I����H.I��#�/��B/��8�^Z�[���r�\��@�6$�t r�/�m��9>�m�lr���-)�i�=�g�vf�%6
#C���Yhb��Zi�r��(ǝ�@8����Fև�J�c ��-gzV��i�Z�:���O�'R��z���0����pcJ�x:fb� d�U�9���Q��S�ݕ��Z�V��(;|�#J�S��n���7\&M�:�S��o��=�y�ʺ��3Mx(`��h=F�(#�})17��^7����7!Wx��F����|��@H�����2��)�zD�N��q���Υ�L���ۉ�L�
�i~XB���;����Ov���^>ӕh*���a�������9��AZ�\П�
����i{�����#;�����pkm��g�P�ڡ!��K���;�����-B�}�̃�L�y�M} �Fu�f 5��Ѯk!��)���Օ5˩�T��x2�^�GC����\3GJﰨ�/�gΎ�u0.3wur	H�:ix��/�J�_Kj��?x�t�\v����@V8/����d��g]����Cf1!�>��0"���~�'+��D3w�U��������8�Pc�����J78��Ƿ�l f;fSN��}�Ԉܫt|�/
�}��D��U�7锬n�(nJ��pr\�Ob��6�=��	!wf�V�p������R�va�͚F�]ݺ��{�#5G���P�X �������(����B���R��9�pn�d�j�6�>~��S�o��M�Ə1�ϯ{I��ʉXn.�{-c2��Ve�q@�4j��v���t�Z���|O�C��FnZ�X�X��h�q��(BS�wh�`��?
�c�[-����_��;[���K�5�x�CO��HB3�|o��[�$T�69���3���6PZJN��\��;�e����p����=t��*�6]�;��3xТ���l!�� �r��5��B�v�Y���ʃL��b��q��]��3�����-Ų��u�6@"1�Ƞ�|�K��j��`H����`����
�_7w8���<g�Ȗ��]����YR��E"��?�m�R�͌,�r
:��nsQ�)����[��E�r8^<;9��nS܉�K�J0�e�Qƻ#]q��ն^s]WA�:̓u�N��6�*�d���ټ�r��J�ӻ�Ƨ���ih�Af\GDSl�W��Ğ�*F+�"Iܐû�<��Sau��`�ŕX�ˠ�R�?|X�XǍ���Y�&q)Y/%��
#�PK������Y�.!�����{�#p��B�����*�l��g������M:� {)�t�6v]�ײ�3BcS��S�:k����W��@�v-/�o�4B�[��l��[��-"�Xb,�9:\nw�ꇑh�!����_��������te���C�V\�E.���-�Eo�X�C������E(�����B��z>->G��ut�hA}�)�;HPP�n���ٲ 3^<�-#1j�"�ΖC�LZ��$�/�C$�������ތO��W��slS�����h{I�r�����C=��"�?��GD�Po�̆JGL�K�(xfh���ܸh0>���8����O��+��N��*���c�K��dL��S���|c�3�N:F��+1�N�߶����:NT[���1P���O�����5���p9�q�Fe��}bh۟��q�H���d����0�PG���T3N��<pP�u.�B��J���'|H���Lɻ�YGܣ�鰅�z��K!	|����]#�F8uc*"��-���{yE!����K\�,���T��!(�M�ܼ�iM����$i��1�!��qҊ�=@ZF������Yn�y��6
#_A���|���A��Z���2��R��N>��H��(��\k+��O��I�2{�Κ��EbUmA����K���Js�bC�"z��,�v�m�$�y.O���5�܃��C×Df���e���6[��� 60vr!�;M�!J�f�W젥��Q��d���h��5�'�G �7 ��4���˶�-Yˍ��i2-�F�R(�T���=s`Igw~YD�@�{a7�~Au����Ia�������1feo-�s�÷]^<"��S.�9Υ��VН�-�i���C��A9Ě?��\����t�Zn��8���̨�b}7���@����#W�8�������*!9h!Kr[ˆ;M'�p�k
�7"�7��g�߭,W� �Fc�:7�s1f���M��߂��7&9���ãe�_�o���H��@�N�A��:�Q�k��*V��B��ɹe{\q���K&�
�D �KfEn-
lv&ܸ��c�d�z�J���p�!Vܣ\y�[߭m8����_v�@A�!7�Q�"�J2mH��Ow���_
��y?�a�˶H eaq���%u�k�y�8��-��l����ۉ�P"�De:�r����Eא��3�f�g*F%�j4��8isL��%&a+m�*�cg�9��Q����j|���m��GI[{2�wfՌ �h�L��n�1����w�K5ُD�+��|3/S���J7�uC��P�i]�^E��LXHS?ˬ)]��X]h\�5�-�ޞ9[t��h���~B��հ��۹-��Q��G��q� ��`���~��LT�I#�X�%���Yg�|ݴx�^��A1oJ���n�I}�S`	G�Ų_��[(P�hOh׎�jWSW���;�2��mF�h���4��Xv������]�BV�V��b�ң�]������x�d�B-�
��=H*܃�0�PĪdÅ�(D�4�F­�bt���g�b�E 7� ��E�l�>�����l�8���ֽj؉>�O��¸g��HiBs�p�a�㞟�������q�.m����Wx��{:0QRk-q�4���cF�c��C`�ڼh�$Q�l��[U��pO�{h=i�����k��=�C��(_�#%�b��&�H��VY�M%�y�,��+f��"�vM`������ϝ�)��Y�Z�m����>q�~�VS�L�lvžh2�(/�3�e7y�]�3(�)%���.$���=��������P��&�8�N�x��>I�F��Ǵ� �)�Ə~�s��^�>���̑�Hq=iS��H�ԛ�8�S^3�t�(���CZ���y�T,��]���ha=��;�I��i�C#4A�������y�UKZl4 ̽&�Lɏ�d��?�)���l�<]��O�����c�#�:W*AcڃXqV-���Ğ�M~�r|�������շ�y���� k6�R�7�]��l�A��o�����>#�O��	�TO����;_eɇ���T��G {[�ĦZ�2ŗ~�7�p�z�\|�2y�8i�����f6#�5�i�Z7τ���dT�a@  ���(��1�/�3�5��"KP���W�����@�M�y��{~(dI�b��Ψ��^�����
R�I�u+(�7�27R$*�&d����}p-x�h�0R�*��r������Cz
�pR�W6�iog�cTtGwʌ�jz"3<�����/s �5E͕jRhY�n6��iD�r��Oj�̫2T���ٻ*��@� ��F��3*I�w��e��_(�1=D�rěW�\ut�����h�Oy/�8�~p^�:�qB��S��|1�f�I���稽�n�HnI�6Q�t�{N��w�B��}}M��Us���@lT9�hD7�E��ژ��C�;�H��]BM9�@��uT��90��7u���Y�#b0�1��a�!��M��,��ER�'��A��7��ȧ����x����QɹĂ��������gmVh5ԝ�v�����%A��L�IS�2��w&�1���/Bp����Z)���,E̻!qJ��v�������-W��,r�h�����3����;�����]H�f���9������p���9��k{b4}j�w�����wA��3�/~�tIi�f�o�r��D���ʉ)��O11��ET���-
S_��t�z��n�ڑL�\f�����ؓcs��t�t��y /zgv��b�Q&!Bc��0W����}�	�����D�<����~��κ��\�x�FX>�V�q�p��m�ļ/z�As����40��"�ۓ��R�"�{�,����$�{DZԕ6_���i�6!e[~F�^[ɟ;2Eo�n}/4 \���qK3�sk��+���S�;e����gb�x�գҝ��m�ݘ���%��#o�(7TAM�IV�i��"$��,k��Z��oc�P6�W��K*����x���@�ĭj��+#	��`��o:�<����<7cb�q�@G&`�6�Q��S*o�4��A2��R�G�9���	��X�8�hw{j��ͭ��2'���ƶ]mWS������~0g~cD��a��]'3��2�'�O��	�D�1��{�'��$��K8���!��`Q�y<��s���)���&���p[�V��m�}���O�I����p*��Tk6glk~S&W���K���h#�e�;?��}^���
y$�: �cN.���s�P҇��<'WX�V�8}��V3b��)�|vN�*KƬ�����(�͘-�)ҏt/t���2\��	��^c���9�N��f��_��U�9�T˨ytB?��LZ<�2�g�FΠ{�����E�h�%R����R�G�t�l龈�[H�V�?_��)�paa��Z^-[�W�}�k|r!qt�|\�<\%c�����~e&q�cݺ��Zb�PK��@�������	���-Lȶ��n����p��2�O�WC����BU<!�����F�����VE���fNv(�EKBIE�a�]�����]���0�:L-���w-Y*�B���,��XDF��P�}-!��4�$�]�w՚R���ѤEj�Ǉjm"���x�2z^:�e|�Ho^_����HKۨ^lP���aR��Aje9R�y�t*.̠M���к�����9�iCdM�����5������PJ����:�A����|H@�x�����ϪC�擌�N��G/+�������\�Vd����_�i�l�N ��Sk��ۏy��$'�J��,µ*~��������.oA^�j�J���t�f(�������z�׍���j����q��|� y�4P��ѸBm�.!����'	�m ���X�<���bt�8E/�D�_訑[�r�&�n�0�y��ay���2��;QAĴ�s�����9pn�3��qZy�+�o��_�6���2S�WF�1�~�����c�4�E'�Oc�a��8b�����Y���L�����EֲWڔ�a]�M�P��������Q���������z���(7�ܳ%�#�b�8���T��`�/�G�vs~;��>Лp���<��,#�w��"�p���C��g��Qye6ua-
G/�����>)���=9D�VARsDճZ/�.�zO��'y� ����3�v��;��a�6�����Y����h0u���,Z���x�yb���S(@r�X���Oz��\E����c).�����K�qt�"���zi[�����8Rכv����4n����^Rd�`b�r����J�����+�CAQ�V�"�tˬ9߅_/*P9u�d1p��9�N쾶Ft&s�A�OBaҧE�\�D�]Sf��9�9�= �~�ė�S�w)�%G��*[�\ί=��R��0C�4�OI�RbK���d �����o�&YJ�ð���W�/+^�u�=q
`7�<��~��C� <�Ea>I��"�_@.FL�)�+bd�
	�c�D����IrzL���sN�����������6�AH�Y�ӽ�u����oW8b~��Zl�+���kij�_,��Vl��R�NܓG�Mea�7'6�z5S���;� ���Buc���[���������;ʛ��w![=P�(���o(�詶m�P��!2�:�����˱�O?M�S��	y-��]m�\c��$��o�HI��CA%��m��{T>�s�GW�vbt ���̄N�?��ɇ#ҵhJ �x������V;��%��f�wܒQ�/ �u�\��H�xD*��w�:ۇ��������3�n�'fʦ��q�,9B�}�j�����'�V���{T�~��N�Օ%W�u��.&e<��������ȃ�j�-Gql��ےw�z������d�n!,�>��/�Anޖ=��"<�|�I��4^�BR��!� �K�u�Њ(a'6m:2/	޻�����ﯦ�/lU9�D�9�(Ն�"H��k= MJ�EQP�
�P� �k��� ��N��N ���?�;����{�c���s͵��3�Zs	�]�&$� ����6�_�5�i��uw`x�������a�ƎP�V�|�F<l�&$��/p����>�����CQ�@��p�w��A�|ne�m�忯�g[k��!=��q����;���_��I�o�����v��`�>��?�&�Mˣ�1�g�h���r��AQ���;�j,q��O&_/�]�J@4�����V ��r�e��	��s�c��T���[�oߙ'rɋ���5���8�G�K����c�Yf�n�+q��=���柛�)�ēyµ1Ĩ{3�������5'��u�F��������A��x;DE0�ҭ'j�1rk,�*�ZS����U��q}��Ż�R*?�^	����*� ��gy��.0_�%�:��v�h��x�)��u�>�mE�*cgO�z�z��x�Wh[�Qk��� ���R�2�b�VP�oD���=��ꩌ�ޭ� ���>�����f\�?UJ���ݴ�&L�[�椂�x@�בZ���|�w?�ۯ?��Bx-�"y�.x�'�&@�$�A�"�9��>?������U�;h�4���0���L��jX�}X��;�G�ɶR�z���20�I:{��ǫ�����|e�8�Ռ�=x9��Ļ1+l! ����ń@�Aɀ�E�y�}��72Q�錞����8p~!���6!g�/�:�����#|{��
����l���C�Ҹ�A
Mc����X�,��d
��|���μ����Q�Q�j�Fx�Q���3?�w�GӉ�&��Ԅ�A�B���F8쾧6WJ�-ϝ1�1��Mz2:�!��sH�O���8~6�1���+)��V�>,\�=��W'�Z%��6��m�Y`	Ke�-�G����K?��Z��G[屶S�jf�i�хk��ps��v���Q8���  )[{b��檔r^�g�D�ʀ�L�郆�GC0N�ŗ���g�5�w��JlC#�Ɣ�|T�C����R뎎T��˻�nay�D*=(���a������#P�מ�S�v��8���3]�/s=m=o�2�:��,�ybv�>8bPq�9,.�	_B	��^���#=�Tu8����N�į��wUT�grf��s\�����_6���u0F
�%�v�;�X�d��sy����������>���ـ��[ɛ��
��L��Kt��<��z��>�0p�7��9v5�y���S��R���Y�2���@���Nv��5ݹ�!W�o��IG�A�-\B�P�~Ȥ�.�7��H�S꠵����el���5UԂ�LKf�����C:DPu&�lk�o��G]g���;:���>�L]��Q�iUY��F�w
���)�_\��̦M�]Lr�\pi����O[H����^m�M9Z��΍ ߇W���=`6��;��\	ݭ�>��\G:��=j��Y���q�N�s�!���Si�+��sb�Z/M�3`?ӞY��	������Ƹڌ2���p(�>�/�`�4y�����k���P����#�Y�!��J���>�zߺv���`W�Y"o�3q/��e��f�v��=Q���[4�Ңs�� ��w;�++����Qn�"��،y���`��F��EΨŇ����s�*�G�6T�0�����L�Ge�*(���R8s��c$���^������b�7������N�mc-"�������H�P-�X}n�I;U���ʅOt�(J���׻�T (5��������0�{%�J�|Zpw$^�aZM��I�������S	\;�)EQO��[���y?{3"��jˇ��1o�ơT�[|jXB�!��I�Ж�0�
��.�"���
L��j����_������Lz�Mf*!v�#͊�R�VB����x��N/�ѢM�L���%8�z�q�`?��EF��qē�[ԫ ������&>��GmB�J�#|0��<�1����aj�A�~]# t����*Ӝ.eh��L�t��C��S�+j���ٵ^?9KY���/�*ScH�<�l�_Z�Iާ��\��$+b��&�O	< d5i�}̫�?��)���H�We0�P��%n�\{��4�7��#@ܘk�'=��[t�mM�]��Q �T&��1f�o2ڳ��q\홭�^3?���6����s��u����R}�7�+L�y�,a�{_q�6�vE�e�)7K��_�4lYn�44B�����Pھk�-&?�>�����Q����Oߐm��x䱈��Os��i٢��Vrs�� �r�1��{�]��͝�!����c�_q"�bA����g�.���(=��6�˼/Z������Ji�|��S9,-�����l:��jm�iT�p0��ӊ�����t����3Y��O��6Vin�3!b�mJ��ѹ��e�ѥ\��2��c������좒Wf����o��:�+����,W���$�]���S��a�z틯����R�E��S=�����Wyiza�s���֨�l%~�Q ��6�3�
G�n�G�b%ݡ�L�̔��|��괠�{y|ħ���dew��J���v&K;�V�EiK�K��j�r#M,�7�B��:+�'���1���m�eK�k�^�9���~r��j'��8ikb`5�-D�sO<�&�9#j�>��k]�!�&t�X�Ntz��x7�_E�qB(���r	�N^���̋�2�oF��ik��OZ�߈K���<���:_RK��� u��_E�Q���j�G^zi�^��p2�:�r������7n�o*	C�Zv�w �30&,'5�H�ni�T��,Z�F�(�GL'Me&#H�g��]f����N����wz��K�����e�dNU���3�@�����	Ȑ�mNR��й��,��u��v�0����>�N]��v�u-�,��W�У�����г^��s�[�v�"�C�G)�5�K��4�����;(gM~�9q՘s����4y��������C���-�ٟ�q�8��a!N�L�@`l�(p��-�O噘��%�l�Z6�(4^��� ���ӣ��Q6.�fi70�Q2Oj_L��[��)�le����������.b.�'PB�T���j���O��J���9M�0go�&��ﵖW:�D���![]��1_U��@C����-�bK͹����T-��dĊ�(�mS|�gENi���*\-jd�bY�H-b@���&���qo�I��lV`XB���M?2t�9��8�Ac�x�C=�����@�K��� ����[f�T���F�O�&�8�0[,��.���
�٘󩀯�e�Z����o�`���������	,krI4>`� 2f��S���C��å�F]o�d�?&2�Ej6"%�ǜ�d̍ウ�6T*��0͕�lV(�^����	*�u��*]w��x�D~] <Qd!�њ�p�����%X]P�o������*x
���l��^�~y�[X��U�yn��|�n���KR#��m�C�k�c�ߠW@�[�fR��Sv>�rs7q�ϝ�Q�����<�� t$d_M�I(�Y;%/b�HQ���>�0.�~�����I�ć`2��b9͵Ȯ8��%��B�WO�ؼl(�D���.T�w���X��|gP0b���3	R̵u�<���xU�gw�5�V���[Q;�_��zjw��W�<vi1[;��]a�To����1���դ
�%T	�������⒃��+�<~��:ڋ'��o�U��;r@7o6W����eYU�%��3���38n���u⵶O�
��B���A��MU���Ъ����B�>AQ�	1N��d�5	W���xW�fgsiܹ䎠ܪ�ڰ�2n�mjX8�T����+f��o�vYv�R�)bQ4f�!D��� �n_%t���)���fbGZ��y�賊-�&���{�bjgP0!��
�^vׁ��Ice�6.G��jO�z�X�&o�.��C��Vز�4�(��4����Jp��D�/g�(�L���ٚ����͛���u�z�H�j4w�	���am=s��Q��NA� �۵ZKph^�������H(������I���|q}�yP[U.�P��r��x���-�Q*Eڸ�qw$w�`�������Q#>���!��_K/^��Y��6�{���2���e��'�\hT�#ՠ� ���H�WKn��߉�f�5���@��W.�������F���4�� ;Ǭ�r�@T����ǫ����~+�,��q���Q�������y�`!�]��R����|	ũ��	�ccPb������0��_,R��HR3�;:M]�
��I��m'�b@�8�g�:ޝB�e��*4��Ak���8�\v\J���l06s�,����v��gR�����Jkm���Q��A�f���lI�!�;1��<}�J��yM�r�=��h7b��5����<�K����p׬q+y���i<�Z�?��$��ڡ�q�qߢ0�N6�%��T�RP��aF+�`mc��)�5×U�����92�Yp_w˷�lsǲU�V��-]�[P_[�*��7���J�Wl!G�k磻蝚h�o�+�\71���k59Cš��C7@\ړ�P�Ԫ|����2
��yn���J�[ӆO+d-w54u�*W�K����@��r�K��l�mg�X;'���~�$5���ң�-��2#)�}��n��e�R�&[v��B!�õl�C��>� I�Z9Q4�L�|?��xC�5��X�4F%1�И��䨆G��Ue���
g�!x�r�AS�y
d՚��d�ZL�� }E(Q�p��K 5����*��L7	J�m��z�O4�� ��)%LqP֏�qI�k��*�g�Koj�n�d�L���c�E8O�)�Cbaf�&��D��5!��3���+-_�}H�^9.�m���P����-�V$A�<S��(��IX��wO) �>:n�w��WE9>���0�����lt��:-�i���;e^m�j]7���%��Ko���7cs��3�k�����Y�~z�L"7�p˰"~H�j�M5����m��E�?������7�}b��<Bl�7 ������qe{�*�S�'�Jtü�q�?�]��#�;,Y�WK-��㹨�Z�:��%P�|W�vܵ��_qjGk�W>,��t��v�H��T�խ��!z	�K
�n�(P}�.���muHB��~I�EbFQFاpkT�ў�{/%��ox�|d4�]v�L�~���km�y{�T��U?�I�_fx?f<cFMԐ�a���V}�ԭ�JP
��L[�p>��*�V�)�/�߳v����z�?J:w��|��Fe@8X������r�N鯵�����&�<�-��%,w!�Pv=}bM�6G��V->��*��=?cg���� �V��$�A��DC����R��eK��w0z^�n	W���޲�>��ڐ����y�㎯�L�⋦՚m�N#��E�}�ݒE3�ͯ�6'w���X�?z4��Y/������'�Dj��**/���x���Ll� J���J�.���0Q:�_�39ǳ�> 9L�.[��O��
�!\���wJZ��I��l+6��KkYsǇ^������
�t2�,��X���~�����Ve�����s�tʅ�l�X Ј��"��r`��O��=���Kt�Ls]H��g	�I�\��j��'&+����Ҍkʱ	j�wi�	��׋�}���*�S���×��Qq�㭊�V��
0�7.ބ�h���E@ ��'itƼA��E`�5�~\�[����X�J����4���(��({וP�;��7F&��(��NA�c�ֹlwO�c|�y9��6Ԇ�GF{�/���.�����-��RE��E��[C,����ސ�]X{-����-�
��	Tn1r"?'oa )26���]���ح�Y��=��Z��7Y�,,��8�qك�O�D�+�ڦ��I/1s��ܼ(�������#�*�0����2�:9n���=BE?+@�ʰ��\�$�h<�0>��@FGn�"��Sc��)��Uh�,hd�M�p̞)H�����گ�M<)�� wj�8�����ɮ���럇ҕ7�*��JG�z�g�mN���V�o VR:�[j�QV9��#�Ŏ���/O�� &G�E�4�Z��j��2�-ۛ�!,����H)�&4���n���h�)Zꌭ
p+��ԾZ�h� ���vv%]�X�W�ں�Ș��5jl��[����\���/D����YDa�mw�"��꼴����J>>GQ��mtD���$I��+���Y�q2̒��e.�υ[�D��	g�^��2�q���&qP� �Z8��*Lg��̶:Ә;ZK�Wv�CV�����sWG�tU���瑪R�=�烻��V���A���7��I����W�[]0&U�w�嬨2b�� �o��GŚ|����o�K�@������|��A��Q�Jܦ�t���;s֗�K�O�1���e+�J�)��H�/ke9���B2������r�͞�X�P�w�}R��)o�;_�_V��4�MU��P�W�\˰V��z%�j�����㭌�6�'5 kgȈ3��AH�4g��(�X��v	��I��t�t�N�c�.\WP���� ����>�$��Ҭ��[Kc��Zq���f%%��� gU����]��K{6�C�\L�� ��$�ـ��Q����Kӵ1�|t��RG��4�Ok��;���&��k��7�k΅���Q
	��h�*\��)�6�2?�k܌�mc��?ޛ�^St�2��c$��6����LM�� �*pj�����J�4Y�k�#�ݐߍ���nc۞��P��j;wh�܈�~��#$��杻���.��v�*9;�4�U�ߗe1pO�����ݖUE����#�
垨g�_c7ܳ̽�
�hh�#��x���>ι�/"��J븕��� 4����b3h�.@x<�[)���**A�ٹ-uՠ@)ާu�k��Q��-Ȉ��l6����ӗr����؂w�ܔ>"�X`䨴�	��2�B<��d�ֿb ͑Ŗ�����Ϟ!,SI�Wyb����Ѡ3J���J��ֿ�4h\��LY��<6�̸�O�����>��m�0aMN�3�$_jj�ܲ%+1�`| A��V7��m1�:7#y_�4�p� Y��ch���+�%�nM��Ծ�җ'�[=�] g!|3h+����D�9F�Qe�)�J$R����Z��v�����v|gB���T*�R}�6l�N�Zޤd[�^��b2#��[����#�<i���_F���g� kO�L�Ӣ֧-�$q�q4ɪ���l��y����^�Z�*@�N��Y�^	7,�;^v?���^�Yb�j>�aH�8�,+�`�ϧ�Gf�H���3C��6�X�����q\�m��i�x���%c��c}$���/�����y�jO�3�LwφD0�R��~���C{�/	Y��2�D��@:��=��w����gMC?��6��:\+���v*&=r������6t=
�.��U�rlNz�킩N������?g�V6� ��)���ݰ:F�R��^���Mj��Y=1�L�ᔮ�P��u��q)LS:��Y���K%�q�(_rI�(����XsԮ�G�Ml���j?��)��T��,�v@&�Ci�	3�Y�{�zUL��kǅZ�4}\�%���@ep�Y�@��NE{�TI�X��d5�1O��;���`�N�c�\��)κ���;�P�@��Ll�^ZTW��kN~�R7�:�fj���q���#�*�)�����j	'��b��y<ǳX��Ķ<9��;w�z�I�G��Mn0�&̜�?��'�sF�Pn�ij�L��~�����mt���'�׹��Nl@XKs:z��jXB�Vv	H�O(�����;\���|�� ����Ow:�YN*-�l�ѻ޳$Lj4��f�)4u.����e�Օ�PvL�x�!f�*��p�S��t*��j{pw��|��Nl��\��q>%n���9���V�͙�4��ϱ�GP��nU��r������r���?�~c>�mC�������AX��͜�K#�l�yMeS-���@��(��|~|���@�q��*p�ʲ�q=�����!:k�
�'GwN�2
�2$<E�=b&>��9D����Dڂ��߈�O�����I�R����ǧ.}9>��ժ�
�z�(���Nz�8������BOJ�~g��� �0tz��ե�K��U�
o��G�:xҟ2٧Ƞ�+��͊���ud�l�]��5hۄ^����u����ӣ�Ϧe�~}���uH��߿����ţ���5�Nl�X|p�ƹ.���o�}����		3Mk���+!�ͧY���<���X���_�?1�SsldЅ���޴�ۑ�$�����
t��Cg�H����-���|���تXʁ�}�Ž��	�R�E�5�)�(c4h7����I%A����L��bb�{5�V��C:�0c˿�C- �fS��]\!W�"�����@���] '�z�Ha�MF�����P�3�Z���>�nKZ���ƶ��%yU�����,~B�Ƹ\�@�4+���G�����v��4p������T����(������g)��*w�嗴ڛ�`�I���"n7-�6����"e@��Lv���P�}��S�f�v����9�jY��+�m5��n+<^�9E}K���E��u��t�',CtWE ��'�n��B��_.�B��ǫ$F�T,3e'���D޳��ߢ���\˚)e��u��03�J:YM:UNţ~c~�9I���*��Hk�#-��M��G��"�!�=V��QȩݴzsHQ�
���vXB�z5�O7K'�G��_�l[�H?��L_��$���~�¹��}U��rn���Z]
[�e>`�9�w��Z�M�@��]0����y��˾Y�Z���!�+��9.J6�qw�ű�'��5�+N$���;��b���ׄ��V��J<�,����c;�������Œ�^eK@s���/><���~�m(�.VD�����{���s�;��w5uM6}�旙W%8Ͻ�a�w���/�"n
�@��:l�d��O�m�]��}�"Ӧe�Ԅ�Ð������~>uU�x��n����4W����{Tkl��nZ��y���[�6Ɍ�
J`����My��k��:���(�jk�S��u_��{��}����;4&1b�oZ�6�\�t��t����'ڴ8G�W�y_
�>��,�7��_l���n!,�`�w����ץX]�XiN	����)��'�+ ��f"W�Ž~�̲��K�
4��9�p�n��zl������s ���Tf_��W������C�&Q�q.�H]��+	��ۙgN��v�%Ʋ$(�Y����k����u$^��[Z�3K8���ר࠰Լ��n�K��� �_�E�?����rG7�[v�s��F��!wu?��hg��fּ�vӟ����hR���׸����J� �s�9�Yv��8e�]8�Mڇ���̡s|\A�Yi'޽^|��~/U�UC#֯���H?
p�~|�2�|S�TK>�P��]�H�(:�X�s�i��K��]�%�N��w������R��߳Ճ��?��S����^�����>u!���z={�^�C���O�av�
�?�ҝh����3h4s8�'���4��Ŀ��B�SGŞ�gH�As��h�ʝ���66�+�<z�����
W����Ϻ���&d���{,���Sz/���h�*G����,�S垱�5T���&}I�d���ob%���t��o����#�y��}��G�D�Bo&��I��ې*)�[CCI�дCa͜�ߡm����y�ۊ����uo�~��r�bM|��-�πؖ�ݴY9:����[ډ��r�o��AZ�6��ʡ}�Fߨ���悂�n��1����G�b4�=�c���RC�aq���-]9h՘�vYK�?N]��&+.SX���n�:���e���Zg�ju����g�͑�\e�P4�VJ���eE�z�Ϟ���v�E�'�2xF*�uh�/������m�&����8���%�9z�ȶ�QB	Z���imwel6�
���!�A/T(�"�o	�k�P��q���4�K�c���?:��o��ؿ�t�{�����n�[[�+���Z+SmC��&r���y�l�jg3��ˮ��ơ�')��8}).�l�`����yK]�s����FƭҀ���®}%F=�u�����\
�x���_#����ɰ?&w���(H	 ��	�-l�	J�Q�������{��
�P��w�)�<�[C@l������	e,��?j��V	D�G7�~���,e+�(ݬ�Qi>m���� t  �g�D'8��@�2�M����YJ�3OG	����c�P�8�����z,�-��8�����U�m�예���o	Y�����w���6�C!�j�Y}>��ɀ�q�ѿ�p.�t+�^����su�=2&n�ي�gé������S�'��u]:��"ms���e��t)U-����{��#T��>.���<������>F��mC;�N;�)�3'&�R�:�c9�\vH�^�SCa�k�	@�7��j����/[��[�����˫z�L��k������e
R�#1�l#�����I[�'��N7���d��lG!���?6�*�0>��!��a	��#�Ujkk�س�. 1czJ�!��r=��.�=�3��m��Sқ�xM�k���&��4+�:S� �oW���/��9�.�7'��Q�͓��P�{ED��z5�K�:[o�ܚ]�{�$�ӵ��N��Y��M|����7կ�3�|{���#`Cu~�)>�駓�[�����	3Ѧ�a���
6�6�4M��!��\�տN��@�:�	����p2C�E�j\�b9���Gx��f��lN"GeH}����*RTw~c"�ti��ཞD�	j�q>m�_[��y�@-$ɠC!2�`_��z`�-��0J�޴h�2�N'f���䉛�K�_� �w��߰�7��-���l���r鯒߯�K�����c���� ���Yi@ۃOc�8��2[_��`w�c�!L�ja���/<�醙��1^R��?�\
�?���Q݅ R�Q:� �� �_���J9t�>��ѵ 3�Vg��*L����
�sD�tnć���{a��W-�lE�[3�F��h��<N�m�?.S��X�����4:�ƣ��5�H/��Κ�n�I�u���Sm{�0�'�O�!�yN�3����NE�l��L������a7���Y�0��2�J��Z����5Ѻ*����04(���?UX�����&��v��N�AZ��4d;"����i�v��7�l1��vSOP����Z�{s�B���Gj�RXT��FDH��I�dq4)�ͽR�����W�K���ܼ=�鈛�|i�cBJ�ޛ^���8֣+�y���EJ����g_F�,P��~���;1bm-�M���� f������1�}�<	�$D1�������M��t���RX�N�]�3�|6�9z�έ~�R���<�=#y����k� �v7��`��X���*bZ�?��6��6�|\����zrΘ��ӎ͔�"f{n�j�X��c?X�S�O������}�
��-���ٱ�9�Jʞcc�� B^&��	�ID�vo
���g�os�5���T�O�C;�,�ߥ�Iig����Z��$�2�I��ҍ����;Ko�=���?]�>�}���V�x�8����M�t�x��$�>�W����I?�m���X�z���d���u�t��m���,�Sez��zp}@���/��mv�)��[ӟ&���	`�Œ" ��)�`/ ��˨�R��>��(�v�DZb��/u����	ѯर<�%���A�9�cG�z�.yŦ�)6&�G�t�'�%�A��� ���k�)�*ʱ��~�O8�$�X� �2�8��P~�R8mS�gF�z~��2��1�ga�U���cD��'�����ȓӈū)��ó�Q��:�+��\��/n�DX�ݲ�|?_'bd�?j
�H���蠋����J�%1,D��%~bػ#G'���]�[;x�B8��RL����]���c�Z+0CO����޼��v���&K\ÂR N���������c�a���A��_�f�ui�~��z|֝2ð3�?���*fS�`�jަ����@R��+�DA�Z*#������k�kɭ�OOL4JR
���.�Sz�|�C��&7uz���z�:}�b��fJ�_�}M��uj�Z�h�4�!�*�4�6�ȃ���B �g��!������5�����g�*)?b�zt蝖��9H=g�Ƿ;ah�v<��2 NQ1/3�2�Hz:��U�f'��EQE&�m`��h��qx��嫦����������gT��=���3�������]i�=�8�Ǆ[��8�j
����əJ�ԝ(�u{r��5�-(RJnzVM�o_k�p�jGv�{����e *i860D��A���_��/�ٰ�r�>D\��j������������͗�����IN�o,���m۝�..^~֌g�o����nɞ�EC�`��^�{���ѣ7�!.�L���ϸ�.!��=����E�Y:	< �_!b���{�-^�������d�p7~���z�[��^i�MQ����$K��s��9YxD��J*֮�,�Mv}=��턈��qsn���Cd�MjLրg�*���Kk�=T�#7B8��!+��5�)x��=9	Ѳѻ��˟�����X���pK���6�S�s#_L��7q�3t���g��yy(2Xܨ�H��9�˜�>W/"�'U6]�@���S���X���=S�����k��;�p1qƗSR����l+��hz�W����d4�ғ�ٞ�ao�� �A�u��i�.���ב{V�xw�fl�L(Fk�B��\S�^Y=�T�t��ny\�pM;��1E�㲯��T��^S�`D��Ͱ3E���@�Z�=1��KƹTi����b���q�	s̡��<
�]�VV�i�=�FYre}�/��(f�Sՙ�;�(��,��]��@�K��,���1�S�5sCU��|�5Թ�vk��w�;J22-zt�#'������aR��e��S[��	i������G��fPs�*7cW��,��*+*���P�q��+}$dn���	�)��s�����@Z=RA�����
��k�=ee��W�`g`�CvT���2�m$#K��}-���� ���l��tS�X�Ձ9X�cX���2�[R׭͋R���na�� ~�aUϜ����a^������܆��W���j�6AuҖ��.؅Q�4����|�V]0�S�bG�d�ȕղa��%�vb����޷FЂ��%�_e��������5ӎ��5�ɀ
+�q�c�qvC-^��&�Y`�sS��t�����z��O��5Zǹ�'�ف����UW��|��N����bgo������J�ý�f�X���eCSVq|�E6����X���(d����xxi䍭�Iu�_��$M+���Q�1�R���}����'�Z�	����<��O��h&_c��7��rA�pb�_OL�å��&��[��o/ X�	��ߜu�m���B�$U�u*}W��MS��!BX��W:��G����*��j�. ~����@AR���o���x�KX�	M�<��(��c�C��y2�}���Q��XF$r�v+:]ɚ�v�M&U)����m	>�ێ=�����/R�-!�r�
{��}�8�����\���s�Ċ�Pw�#X9��������
~Uu�ܘ��@���;j�~�L��~���8��<1	Z 4V�A4�7�#�nT.���光�����C�����(��X�i�F@��n�7��l'�S:N��k4@���?����M��nR�gM&��I=1�T_~�-s�����v�D���+�(�h�\M�Y��U�6ٗ1.���naf�O����=����N���*�!@رF����������rW}aܥ��B�	3RG�f
�?+B�b�*�sC�s���8o���EIԻ0Z���9�28)+=�e3��h9+���0��y�]R��@,����ܤ�(K��4� ������\Y3���~Ý_ľ��/z"0G(��A����U���W�i���H�esx�O���X����8&$���s}k����ykY��X�ۅ�y��h� �蹭�4�A/���c$�]�O���/=�8Ӳ��t!눪�F�8W��~�U{=JZ��l��f�-ԏ=�������K�Y��d5�tz?|[��F���;��2{��9��倨��c���:����xLl"C��A��u\�s*u�� ��d���v��U�W*�\�‖aNm�w``y�{��9�j=�V�Y�����1�lu^6��LԌq�k�"�*rR	����u+���ǆ�xL��F�v���a�y�͜*{���%�Z3�rY�AnT�S&;�j��/*1��]�&�E�9�}p{Ԡ�cw#c\:\��C�!�TڦH��uv�É|���x���a��� �n_p.2�+D�[�(����68湞yT�a�:��Z�Mm(E��n��[�ٵ(����T;��lbz�3�\;}D�0��%��}�B˜�E/quL���O����je�~c�W`yf�b�kR�'p�cx�+��?ܵ����
�g�c
L�u�Z�e��m�`gB
gM���) )��pBFW2�qD��B���1�-�_��}!A;b<=!��n�o��?B�6�QZY� e%d�x�gE��X�Ͻ�Q���b~����֍�x�ج/��^fW��"���s����d�wɩz��1w��=�o�^�Og��k'2#���Tʱ�!�^�q����/�0�(��!3��x��m�J x]\��x��;�qLM�Jx��[�%�t�ꐷ&3�iy��������c��/g�L!�*�HayC�'A*H̬���r�7�O��E{��2^�!�a� �5C�S�+�aK�����`EO&߰��F[�kM\@��HM2�T���[�Z|;������,�q�@  PM f]R^/�z��(����uyU]������~��e�V�y@7�?�Ԙt���M�Ll���ƴ��m�se{�<��^�#���%�k�U�����Վ����ٳ�U��������YZ;�mm!����	����$S�����f�1�[�mm`�KD��wb���Qt�e��΂ +5�j[v�l�[���Vsc3o�kش���D�n���g�W<Q,�b8��)C!�.L�"��z����6.P7�܍6��&�vD�CVQ�k��X�(����ǲ���Жd��s�q�ILْ�/�2*��#cބ��7��]�[��W�&\���P&� ��/`#ea[��GC�6$���/���'���h��{;�i�k���/3���b��j��Qs��dP<`P|c�� ��7��@H-}�Q5wAe%�%����7���O�n͒�>�?J�[P�)$��aU�1�}�)��=����h�cPc�u+�:�[�a�b�j
��W��EV"2�V���y[�0�&�i6\�ʍ��3o�����ّ��U|0�]�����$��ZF�<q?Z 6��i$U�(kA����`'�%jV�_�yA_��ٯ �SX.PݩD��/$a��b->H>������Fr����B�`l�Oh�wx�T�o�^T�Ii̻��E=���]�%Š4e�igl�(��f��a�K�g>����_�j4��l�w�ݱ�o^^G����ܳ�&���)�^I���Ď&6�c��J�蛤=��Y-�x�@�s
�DCڰ�
t�����+��r�q�"��`��ϧ�Y)����J�f��nU���$���k kz�m����)������)+�:�L���[�OR!|���I�y>�n�����r	"oA�
g�X6���>��ӦE��W�{:�C�o+�t�"��CL<�z��>=���R"�w	 �����O�g��s������Jz�Sv����b�d��k\E���R[';�|>���U��G쪕BU����	�9 C��ga�q;�h��`?S@e$�!VꞄǭ,i����y���qq坝ܭ�6f�yo��u��eU��ߘ)�m�U�K�kB&ߕG��Q��K*g�D��C1��?��VF������1���֩�E��8�� ���X��YY#�xoy�a<'��T=���l��F�dEPt�����E���,�m>/��"�}��䄇҃K�כ�Ӡ}��rM"4�s5�®x�V�5h�����P?��SZ�SFҫ�P:��Uߕ���H8B*S�����є,;^����A�n�;��m���0!��E�)Os�ˠ6�0���z4Sk�wݤ���;�&#������ʿ�MO@"�X�i�u������ķ��D%bً�Ὺ�@c���K��,��$Xx�=?��绶�(?����H�S�&���Q
�gA�ף8
�<�i
4��`s�
Q�J��%]nu.#�4�����օ&3,�P*�17O�W�i�:J��CUN	NH�{޻��c
���I�&3��f4�%��f5h��Z�1����0��P��^���q����^�����=��Բ_|�{�&���5'�Qe��a��B+�6��&$�� ]�]�t�|[��]��zʬ��J�l�`��N���4Gll�d��%�����7�T1r�eן�oW��Z%mqs�J�	�@q�'��J��#�Y'�F���ĎӾ�n`�3<S��m���7�nG/Ր�2Ӻ�T%WX�ܑ�}�ʶ�4���c7����G�%&|t�4��]����o��I�U����ԳO'$�+�aў$_X��َ��k^^�4����=S"s�+����-����⩨�& b-K����?�m��}s��{Ign5[X��$��J�gU9�+�
��~]9�|��խ
��	jf��)2�w�5�;��jZ�/u�:8���}�wdɃ%��Kː�����m2��j:E��δ#M��@ έX;?ύ𱺣r�ϕ�nKYd���ڲo%�XI�H�~<޶�f���i��Hf/��3y���x��3E��Y��7��������N[�}�QL���:.��}��@k�,�A�FED:����nd�!9�J7H1�H7C�4C#�C��P����}����׺ם׽��׮�[�o��b*p��B��s\?2�]�'�d\�d�#�4��o Q����V��~V<��e���!�;�m��?��Y���A��f��ne~Yx�2t����M[�kƁ���]� ��K�Rl7/����'�_�8��v��W�'  8��+!N�}r[!��]��?"���RM���7ɛ��	ː��_6A�@t��Zxp�<OL�Nj?Jp��`��]%D���8��U��1�(�4�r��]��ty�P�h����2���u�nn@@2F���~j�b�g~��(��9(lϭ���j��Qo��X�bK� ��}�w�t�`C�4��p��Fxz�Gfd��ps�E�dq�$Y�&*~�ے�C��3��:�p��f��ea��&!�XQm�޻( *GlXBDEGW@'{K�}�FDog�ac�ߪ�S�5�s�e3V��2f~=��YBN�� 2�����a�u֊�d�/��[��rK�ŋs��/�p��Z*�en1y
r(>��F��Ab��Π*��wBݛ�B����>�oo]k�޻�	��P�o;�3�A�����R�¶��ϤHߋ�&��ޯYJ�����W�hH_��e��:(!��E�Z�2��Ea��>���1�FW�#��X7͛�J{�o�G�:����u�8��1�j���K?����UU[䥟!R��΀avÞ�x��~�M-n�*#g�fM�� }4`5ϧS�c�c<
�J�'\g�G�j��4�C��/�a~��x�ˎ�7:2���[��7��V��¤��醈�
Bb,v�-�N��M����y{�����9�{�1H�������=WK)wJ�Dl�]�4��I�~�/[y�,ƻ�;��@���j���q ��N��6ftS�P�}p���u�FL����
������z,;dY~��X�@[RjU���i�TQI�o��N�;�������n�bDZ>\t�p��AV7��*��K��9��W�v�WHinU@�'�)��9ׅ�ac�a)��ܴ�,>�_����Qai�I
�x�1ܐ�Q����cw�ʬ�;�	�7��ȪG,� ����7����C���B-�4�5�[��bae�L� V-�#r��u�/	���T���f�8�v���n�u�9d�_���{��ټï>��6��t6�(��l�v׎Y9gA�_��O��Z����T��bǗR����S~jW��C�x���o{	��<�B�@����Z'�D����l�������Sp�q��qHt���i6���W��u��D6H�¡�L؇a�$u�s�0�J�ԅ�=ׯ@��ZkNp���a���h8[��+h�u���O�_� %\!J��\��׫'�QiN��v�*s`k㐫�TeԎ�n+|*e-[4��d�t_U�wU���5�Yv�b��+��s5��(�lq;�04, S�����6���k�������c�^�v�a:d�{�W�:��§��3sJ$��O/h�Bnd��o@~/*e�f��V�X��{2��Ŭ�͗�͘�{X�KH������1B�?�?>H3�����;��z��O
��Iu����N�00����2�P'Kú��3�p,�)<>�Er��{?w��B� Nb��ydl�Yu�� �_\?��7:^a�n�Ct��*ߢ�`�qԄ5�v�Z�#�T��
�?�7)Q<�Ĩ�Q�ίT��n�Θn�gn��/�$vN��N,��U�V�1]E;E�L�v�I����>�V�qku�5�z�J Y8���Ac��J��c3�]>�b��[DL� h�BWo I�h�1�A7S�ET<4ߚ�(Ѧ�f�k�-b,+|q��F2���Ƶ��t*�N#n��,0�	ȝzU��t�;�fT�噓���T����Z�mw�]!�?���J�t�+��z7a�B��w��
��/8U<��\�I��_�7����6n]՝1���t�4�k�0 LeԂܩ�kO�I\�fY�$=4�9����m�f�nD����\TG��昵ނ6��;Lq�b$��翫���.��UL���*�Mrd���ڑ��	bͭY"�rX>&����UL��=u+����_��6n����[)�B��o`��1���!}B>�x�&(6�ãtL����ufP�n���}W����,Z�&eˎ�X�;�i�}�Fb3��1��u�gE7J۾"�|x{ �߳jtޔ�n�O�զ1T8�
��,��K�jK���u���n*��#���a������.Й��_����o}�!����됓x$�fYo�m�0�����dM����`h0:�,B|=#?P�wW��Jd�,f/��[
5UҌ�.��؁��e�*�SK�V�s�Ahμ�j1���]�SQA]�� 9aX���;X��wg��<���������߈v��z��٫|�P�휉������N�?	�������3K)fw��8����V|�ZP��:P]�1�÷x�&�ʨ�%
����l��2�����@D׃�u;ߊ���;f��������[;&N}�I�Im�;
�I���}���QIh*��\[(�XPg���1�����'�n�ח1H�F2�$]�ڱH����n4�?.�s���	�[2��v�M��E#��7h��^ݝp��d���S��yo܈���z�q�B3�U���^��L�a��k�b�8��Ҽ���#�Qx�G�/5��]=�)Е���)��;aߓSL��9>PA��&� ]�1��݋I�ٟ֖� )~ub�[ry0y����VL���z�D[cPXᚥ�K}�����<q��^��n�+:�C��z���U{ٳ��C��w�V#��Mؚ�]����זj	ji$�u��o�kK}"���6�� ?I�_�y$[d�\b�ii�pl�|s�"��@!�M�}�D�|]`���Kۈ������`�Q����.�" �����R��~*���`�R�Ua�D�,K~Q�e�����%��p�:���	�B�Ƃ�� ,��K�[��.M��U57�6q��1�����A�ak4(a�nd�����l�<c |j�WM�I����G��J���w����&����� (��DfNyIz5�L�[ԍ��'d4�?2|��T�
~��-V�T�1ӣ��ӑC(�[���04��C��y��Z3B*r;��l:3+�3�O�>�����#	݉H�D���MՋ%5�o��,�I��� d�^�/mj��xaDh�ӸS[sm
z�֝g+�{�U��P:�j�	�}b��[��X�Ќ���l�l��e��d���;�o�u�CT�-�5�r��@��6j�K\Z�񿴩�#��f�jC;��y?�]S��r��G١��7�y Xtbh4��=a�q)��t<%1Y{),���yrxN�6��sb��q��3��n��5~d��7J}��BZ`�*�)uh���g��8��:X9$�v��1��t�C�5tN�G�}��fiK�uwy�Y���~��/͓�uR�?M֜DØ�� ɷ�gk�ق9��N����X� �舃��2=��'�PE-!S�ŸKcs7omt�r�9���@N�A��,���c��֐:�U]�V�����%�K���E��j*�����Z�'�C��{�Vbq��i�8��6;T�ܖ���1�����]װ�����S�,Õ��0Wr�n]�X^��)�c�i�ۡ�s����RU:��NS��O�� ��^%�]׽NMIw�{˷�?v��!���В�B�.�d�B�����T��Zə�8R�UѤd}8g��賷jG����rzE7�)���׼�iH���o�]�l��]��v�f;��VT���6mZv�y�v�:p��J����e�4WP�xb2�q����D�����Th�`a���G�����$L����4Y��/���"26[��겿�C�:�Ԙw�z"��(���V������t۽��=Y;��m�� ����y>hST�z�O��H������qE��T�Pq���-��H�H	��Wm�D�k��R�aa@���t�zm�'�K7f��{Wܡ�B˩jU�\�97k���2�9/�Ɂ�����
��}:A}=BG_�l����n��n�Ssh�|vd�����3����g75����ǰn�;5��@�h����_�T�S��*�4�Gn�펏��,�|C���"���i
Nb�<�7�'F�-�����Z�����t����P�o��?Rm{�� ���[�_�m`�B[H}�,��_�����~S�[y��%��!�g����4�	��	��w��qD���ZFC�0��Q���E�-o��2V� �v=��}P���
R�K�F��( /Ց�uv��FwqL���.�$b�]3L~�d�je��=w�#7c�0��n��@�=�>e>Mi����m�i���٥�X[�	����-�\�;h��Y
���ʮX�)T�A�߁��{�w���F�����*�&��;f]ֻᆧ.���c�yM��V�ݡK����3[8A`�y��u��y��j�/ڷ��0[��U9��vI(#�,k��b�ƈ�Q�ӊ�ޔ�!��
�p����js4C�ߝ��������YaktT�E�b^أ��/m�cb�-�.�hF.� ��Y�����f8��HK�gҜ_�o������F��`�媒�>!�����]\�2�CF��YG�{��mɢ0�ٞ�J��/�߻��'�&�r�.0��I�s��`�n��p1j���B����}���W���x"�^,�s������a%���7�Q�>����3ht:qE�"#��Ƹ�vV'��,�q<
][Y�=�|v巖��E=GFԤH�d�Q�*�L���j��:6!��#t�훉�۷�7[��vr�$ǰb��}��J8�@�G������C�CM@�H�6(VA�eOZ���1�Ȩ�<h�|�6$MLN�lS��UgT����懖Y̜�q�Xok���i LL��H��kw�,��-��f%g_�Ifb���"�����X�� 슃.��X��g��|����Xd�'�$?�_7��I;�m������=�҅z'?a�@�q�������8a�2�ҲY3K0�3��OM/�A����߫Bx_U�Dbc������U'P�����>��@K���g�5;s`:��q\�5�֐Š��p����:1�Y�p�x�� `��>]!���J����!���ꫂr�e��Usڗ��n���7���+f�/����bOIm��`�G4��s�z�1�Qs��zh�?�9�������ͪ��>	�z��ܷ�7�`
�qu�D� �F~��rYp����3d�S'f�]��m�=Z��D&Ğ����{lv�6�z�$���e6o����;�hJc�~��{��J\�Rvjό�2j�ބ����	�؋��[=O���0J�="�r�W��}k@']5�m!��X��N���3�,97��	����r���	����%o�3#���}�l�Ü���H�_��a���j+{� ������S#�B+>�~��<BW��{Xǧ)��h���������v�}yl�����"�~�u`@<���`s]\+����q�{��04q��ug@a=,<&�S�*½7�a���������� �-P�j-!��Q��56{�����J�.�ƴ�3_E�W���m^Y_��P�SR��6��h�z0Q���R��"�����m#��]�g��R�*��U
HU����A�JA��$���E�Tm��,����P+[m���M'a;�cL�D���U�Z��%+�_��-��mhK��2]���C�ݵ`���F:�_���+�D}.�4���eV�SA�����yX���H��ַ>5��[^vШ�?A���-��AL.��69̮Զ��P`�&�4a$�>���p	��	�TL��Mg.1T��l?&�T��h��^A��&YU�:��sZ;����w�+
������l�a������t_x�S���*�3���R��A�F������C-7�R9��7�Z�LuF8p	�� ����Ԇ���|�!���+v@ya�.%iJ� ӌ�'t��g�_P���R2���p�����-��@M�D�3���==U)��uĮBC#��~=n�w��Ue��h:���k>�QKg���w���Ah�!pd����;�f�_�i�lUi|��m���1}�h��+1�%�!���{_n�«b��!�J7�`
r�<)�����\.�j�K7V��2������T�Am:Ƞ
g�r� ���7���d�Y6X{���(1Y�8�ݩv��_k��H�&����6�Հ������V�4	@7��x���eC9�^���y�l�KMk%*�c�i:�7t���{8�pyk;��f�r�z>�y��?I�]hf풊��i��9�9MG>dpN���si}�\��<i���W�����G��(}��&z��b����& lKy�Bjl/w����SU�+�܇7�X���c������P��Z��HT�:Ú!C���
�VPn*�\aVY��kCᜑbÞN�w��5ȍ�ۖ��>p��0� z��c�ϱ.���r�k'�%qo����B<l��k�x�g+����t�Q��u|���2<M_ҌM:�Ĳ<�LZW�F�P���nz���_I
����/����^�� >}2^:N�Ƚ �r&�\D#ٷ	�}v!C|�(^?ROq}�`a� ,�*���ZLp�$K�p�HQ�Y���[�\�n��׏d�#>�F��~|Z��_ݟ?�Q-K�Ռ��.�e�Z�T@��)��b����j^v���M��D(�3���,_	���0�����2���Z�
IA�i�&��[ 
�bzarzm���L[!D_޸�: _9�7D\��	7o�ji�l��@[��Y,�K[�Y@�q�2sp.Ԧ^�\;R	����Azx�a�����Z�.Á_'�����M���T�$�+�3Q�1���x���YH���eF`E��ovk���f�3khi��=v���u t65�~�F���5m��Y1�uo&�i(�W
jo���t�΢����` r�T;�A,�I��[�E��Ƙ!�$@x�f���*�p�e�j�3�i+�^����)��?�Bh�m�Trig��y9�g����D�hq�@Fo�/��0��ȕj�o�]��Ƌo�v+����]�0�uL֛�d���!U��բ����5��eZUQK��F�k7�0a)
l��ٍJ�o�|�y�@���E�_��9��w���e<�*���qv��#�{P�<����l�A�&PJ\�����v=�k�"��%��Y�\9��3j*źL�٘*�.�5|^[��;���>R<f �/�/��,q�[������;!�}3Z�����Cg�⾙/c4,Ef/�9�J�Z�K������Ӆ�;�c���_��`���/��3�q7�:�&���v��Z)q�q.�&���<����h��K��.���Hv�o�.0x'Q��sD��:�=���0�~�� ॎ���+&���1Q�S�;8��8��DUܘ�p	:�c���>�P5�M-X�Shx��QUf4Ptm4���h�w�'�����\���a���C�Zm��y^{�?�k�+��؆�2�r��0�~k���x�5�W,����ˆl���
-�_f��d�탾�C[Wӵ1wD�>�}�:.^lj��C:�/�����{���(f`��e�����xv��MgwR��m+� L�`���ح�f}�E���+�A�B�G�O���w�]�Q���ք
:�?��m
y|v�.���-soL��?��ݏ���@���b��&-"L�]p.伏!`�7a-�h?�e=fa��psVS��m�H���aVݲ|�z_�[5X3iZHz߲i뚆����&������ˉ���.rcb�@G��x8	�9�ʽS�`�S���=�e��km����m_�����*w��Q��p��)T��ToR�>�����2F퐛0�e�k�G%l���JI-��L�ſ\��t�,��V��鴿��9gƕ��x-Ԥy��-t������Ztqq"^>}�a�����[�c���U=�[��x�v���nbr����-��)6n�F�&� �6��Ê�sY>�/���q�z�,�r�Y���=���������O���<�;�J�N�@��	x)�s�^���%�q���v�7")��{��r�zWm�r���x�������_�Ǉy���ڃ�c�(�B�5����>���ٟ����K���p`���TR����J��� P8�MLT�����۝O��+HIN�?���a1�$c3�%��(�c���暒x:+f�3��[�|& Jl�j]��t�����s7�����ƃ��ݷ>=�&�_S�/��+5����DU�)J7b�kׂ�� �ub؄���F��Dk�x%x�L
;�Duc��T֧h2ٚ���a��"Tr�I#����bNDO���B�1Eo�ÄʽK!���C!5'c����y�"s��~˟����O�m⚉x+��Q�H@���˖�ӏK/�����������W�ol.�ے�1��h'�љ;�U�c���4����S��&��<xy�Ҿv۟m]�!I2������H�Af�V�5���X�,|o5�J���Z�^h��^T�j��~���
��=�b�B����i'l� �a�����b�_�z���a����D�W%�׎B����Iě�Þ-��������+�Si��{�g��;QJ��$X�_W"����W��T�%�dw�zq}���(�궩����>ZMa�|�Kk#��[�n�%ˡ�)|6�X�ƃ�X�3�iƖ_��\և��~Bw�ǻcޓ�Z$b�*�*���N�T��4���2��p��yz������̱3_v]���만y�ca���a�����]�=����[n�4�]��s��#��Ae��������v�a�B�����J��p�G!jCՍQ��V�����q(+DF�ή�ds2���g�Dz�Y�ךb��m�����N������n�z�ɍ[���'���;?� ׅ�˻�VH��\\M/��1��u��A{�m����H���@,��:Đ��&�=�^ʟ�l��b���K,D?��W�nF	ܸE�ٵ���.�a�PfvwR���������؁��@�6��**p嘥V�&.����l�~�'��WQnc�.G;���#v#o3$[a%�"�<�1���0/���S�\^�#j���x:ڨ�	��t�)e*�\",v85W�F
ĐǍ��w�˯�BIr�S�����m��}����B��}m:݂2��./�Ì{�Xz:�]�.&�肐m.?��M�	j����-,i�؀��W���d�?8�n����K�=(v�4�a������6�v����K~�����̰M�Ċ�M$���a6������G�N�eN�c���[��UXV"������Ԝ��W�^rk�*���U	����_k��Ԓ�%Oъ9N"�O�a������{2nc"����L�%G�
Q�-T�M��:�ԡ9U�Ǵ~�J>��#-F
��O+��ҰU����hgs!��VE�-��f����Oz�M��`�x��Џ��0형��9زs�^����q������aW�>W7�O�k�Wȴ,p8��/s[��F�O�3[OtV�Rk�?s���4���B��=s7/�L���������F�/Ϧ���y���L? �L�.YVbe{xJF�	�vZ�S^1�^�Ԃ��<��`b�!&�����VkAl���]~�h���1>Z}y���D��o0{N��9	��<�Ex#z��u�x�t�]��'�^Wم�tr�%�%sT@y��h�ة|[.+�b��Z���J�����xz�~:��:i���}��p�L���C�u�
���]ƕ�C����.՝��a=�%-�9]�1�F�������,N�nj������VK _���q��vZ=u�|n9�f�U���I'�(%\d��Ϗޭ�\��\Z��ڒ�ľW�͌����6�V��?Q�~g"d^P�q���O���!~ 0����؅x�\݃JQ:���y�?6��Q�ˌ�*�_D�&s�j�!4��}0�� ���n�}/,O�����tʷ�'2�נ9,�ݩ ���Zk� ��THX9sҫ�Q�<n��,�V�};��v�5��Uj����ƅS�s��l�� ���n�����F�˖��5O����m�\dۅ�w�A)B��l�t����DP�F�~)�e9��E�q���7��������������2����4�홖�Z��?�����dm��<�	�fd	n!�0�@mG���!�!,��Sҥ*�_$%&^�>�����
?	�c6��X/�N�^��AlY�����b3��T�C���Z�B*� 5��2W'��6��|�sz���ӛf�������OfBD�^Y
ŉ����PsWZ�p�m^��7��=T���D���X�4	��_�/�U@���|Ǒ��+Yu�f2M2H�ы~X����Q4����{�'�V6b��؍)�����x"O���F��0X���~7И�v7�s�>�������x����!�*�i������ܯ�i\�Ŧ`g"�ǭ�����C��z�l:qn����	/���􊡎��bgO\�5�@��p�#�R�<݅�z#�7��N:�'[�+aV0�fj<gpˇ!ryo���߫�=�
�zw�)�3@��Uϡ�x%Oh�����Y�*E���/�3O�N�*�/88�%t�����/�
� O!����²��T�[3�� ��/$��_��1����5�`�|�<?|y��z۬��[�	�U�@�Ъ���>�2����P����(�?��`֤�vk�L�~��Wآ���	R��&�i��R��Pi��^{�3\wk�sn�NW��D"�X��O�u#F�>3�@B��:�
�9Év_PU��*r���⎃-Y�����+�.����T�uT?��_���+z��C����31��zr*c-s��{�t���/�=a��P]C�Ջ��v��+eL�b���U�~��'�î�D�.F�EXuv_�VS~�}�a٪'�:_�e�I�/"G���f��]J"�7s�P�EVꜿ�Y�أ�M��O͋���A(�����3�d8��.��Z&J�,�z��p�EȮ���s��)HY����l���sD���E����9L��0�+@:x��3������!�g�9�g�Ť�p���n�m�X��Ww�;D�tKQ��*K�����:�Ļ�A�߁��D^2.�,����G]��`fB'Y��1�YƯ��g�^aיv�4O;ս�v�z�P��or7��.�к�·��^��}O��i���K�.[_ѥ5��/G��D�_�V��+o�c��|�`^/���#|�T+����^�׬������M��]���dS
��rF��fu���+#5�fJmN��]%���h��&1�N^s˻[����Ò:���ӧ���̀	�����"cO�Ny��-�kU��n唐F]���\st��g)�$��w�l�չlR�?����Z�D'bU�x0F��L��e��HI��#i ����(��@^ɦ�H, �!V=Qz�����xm
��
���OHû��s��@l	+�d��u���N6N��M�aT����S��֟+��	�n�'�Ph'L7�D����C�c����r�Y��d,9�b��4p��S��f�4�l�Z�ZS������Sm��2��2�|�*��Ȥh60�&��ڮ"�-F &0"��K�f�s��*<bh�r��'�B���M�~`�ܾ�h{��)�;�C<}������]]]ŷ�wug�3t��=�}���#`<��~��2O�v�1����-|�՗���&�7?�!A�?�G�5O�7���Z�knfff�V��ӵ�:###`)��@���/�H��ԻĬ��,5�=��1{��[��812Pf^�Ք}�̍�Bj�i�.�� f��*����w{������5*E���Y%f͘X̫�Aފ��׆��>�|�h���dӛ1�b�)<���Σ�/{<Gkd�/Xf��-�&��?#UQ@|�h�Z�.���0j��H����|���p���l[ݔ��JKG���C�������#�O��@�4"�x,��αz�Tnp�(!�2�>u��=/]�/��UǨ+N�]P��|�����@' �����g�	�-\��*�X����K �Oӑ�����<�p���7�u�e�!/73�ۭ�!�m�=,�1�e�z[寵�?r��2W-T��L�����gB]W0n)�K�\����Sg>׽spt��?A�L�3n|ډ9�i�6$���ķY���}�y�j��r��Q�(y�T}�|�!m@�wF&�"VN�QDH���Pу�
��8�0(o�
;yQb�@p�L�lX�Bs�s/F��v���⢺�]~1��� �v�KD�l�6Bh�u���kн��8�y<|�>��u��6�o:��j<k�ER������}�c�`J�JD�����T�`�۾p��/\��.p�0�|��Uڣ�����P��K9܋d�8��Ȱ�f�!��`0����ޥz�Y����oJ�J��#9��X���ʂcG��X����>(C��N���u���@�����c�\��#Y�������4 ��.�����(Nb22��g2x�0���U---�w@1�o�3lo���B���2��ejjl�y�������g��PSS��Y?~a`����I�e=�??>jyu�����i�������������e�-W=Z�G�Qw�}�H�R���'b'�e��	/���rA;�����+ːZY9NU��!q�xȗ~|�D������0: ����=��sr��+��	O+������߯���yt��M�G�їN�=6���ܮ���3_We��z%�Խ#���l��f�À9�:��fgRg:���U ����xr������c=�[{o��Z����Hn�f�2 ~ߦ=��Ë'�/xo��Ł@�7�e4S.�#�?�G��,X���?uL[��L@��FCЄ~�&~ �$���x���s�����8��QN_���epx8\�"��" ��5\��0 �Rk���u`|��Gc�?8�^~~>�x�P ��s��ŐlZ7�g������vT��R�6 8�\���ޞ�R{QY��C3?�0�q���?�145m]g���p�9N���� �b?��.@^I	P��5�q������<@�����p��PP<A�)�{X]��]3>�{{Ռ���r�����u�]zpw�?��^��D^AA�D��+џ���&��s!�{��*�-���a�;���k�@��KHp5�����/n��4*:����G�RN�^~F��s��Lv42}�2��~ ��͏o�I�u�z&�ɣE>���7�t���Ŭcu����؉���7_��4����ϕ�o35Ǌ�;&�(���z\��>��t~����hi8An����GN	���1_;�ҫ�e����U�<�)��})�G	��[�3�	QQ����k��b��>�@��R0���a�jcԶ�aL��L`h�T�_��wc�����;Ƈ^���|S�}Sy|Q�������)Wq�k�C�bN �F�V����w���B �����JO�ڇ{��|������|�*�ʘϴ���rP��i�?�T``1����*��#ӫؖ�����L ������xb����2%�+*^�v�Lu�@;�_�pP߆�$}��@�Ƶ�!�^�,�!�r�P�^	�#(���8�����1�3�!KA��=>���TTll�d��!���������
Ll��96�8���$�һ��d%���R!o�Da���^�4��U���������;0`��/�]>��7ܛ���msl�20y�co;% �h��=��I}*|�
���(��_�\���vѢx�� }�!��i*��7i�3���7�ԅ(��w>�\�*f��H��d+e��8���P�3���C�A�<��:ٹ��r����n�99��58����?d�5�;�����$��4U�J[fkM<�QQ<b�p`(gϿ���i�y�S<���u���,��%Zy�̌�*�51_re8D������۵�~�{ur�ϔH�C|�����"�ҡ�hCaˋ!1@3h:f \��,(���N,3*�O(ษݥg;`1�V��-����֌L��q0���f_
�_�M�<.�J'���L�� w����| \ؽD��Gk ��8 kx^���S�+��@�O��k�������v\�oZ:��Y�Td�
�4�,r�C���0nF�r}u|�l͈�ݖ��.E��2=��0�4���Z1����Wyd����eA[�()���-'�����9Bg�s0�g�u~�r�7]@�!�:� �9F�Ϝ[�nb�Ӷ���!��
J���Q�_� y����B7�`�@��ث�`
�����tQST����y�����g٧�����K��30l��?�O�3G]��,t��;=ج�u�ju�O���D�S�Jh#�v�#
�fߖ&�Y0à z��9��E�p���W���KT�)�u���S�ĝ_���I���ԗ.��?�	��=%e͕|`���������{���䩖rpa~���#
^XZ�Њ�L��'���%�3�d�r
�O�+(y�`0� 8a߇��*d��
Dd ,�^�zTu�%p��M2k�lFښ�Qn^�\ǧ�R����p��p{��%�������)��Ɩ��SSS tn)����A�P��`>��J������s|2؊L>ʔX�?�g���6��q͗I���jj����$��8(��t�̼L�r����.��&�N]����i��h���mT�I
�K� ,S^S�� $�{o�v�	Պ�XNr̒⟛��J�NڞL��@a_z�%vJ���"���@֫����'��㝪�F ����G[��Q�w�~Ei�.p�ʌ��;��i[!:a�F��L҉�F�U���J"9#��2��cY
1� [3��?��Q[�����Og�dm,���Y��((��0I�-�qI©�<{�W�p�s��n���a~/��~�}��_�5��/�Cq1�i�Ƈp+g����i؍4"l=����ݻ�Ʉ+���`o�톹�[�j��`�e�1��F�<�#��{�Q�B�S9��V���\��p��/g�ytjf�(V�u����<���$�����k\�z�l��KP��Ӌ\���Q�T�*�
������).�[�}#?`��*�����J�
����Vv��(���B|����I'�x{:͸T2Q����=������ʠ�w�]Ļ-��|	�bu|��Z���y(^���e*�~�Y�� �+��v �ƻ�A��P;��}�M��XZt`P<���gݹ�#+�1���Vej�R@�Oy���=c���9��\�2�AE�Y��gX/�9X}�n1������\pv�@��{C�O�:i���@��{ݟ��ƣ7��q�Bd=�Лz�Z�|-�ym�M�r����rJ����+Q�L�	I��s0�	_g�DODT�G
�<�Z8{����n��ľ������Mn��^u�(�g'D��7����	|G�V3������zY�C��T�`.��-0��X��x���63��v�L�q�v��Y!ΰ��X����ǰ��z��AV'4L��PL=+�q���Scz��_	��~��=	Dnf�[�z
d:%�°;�Ղy�i�6oE�ȿ����l)��aW�xz��rMJ���)��W���F�wO��&^c6���Q��xF�N�o�z�������!¤
t��k� HO
�(��Y0y�甡���:H|��2�0?)��Z<Ӂw �i���N�r`5�W�$�Tk���}XY(�q�?���"�
��А:K���7I��ۭc�Q��H�p����_b�:0��%4�)G'N17v������>~<F�|�ȶ��JB�^\��,D��f�b�O d�tK�@�qt���$xM1k�c��~��ߤe�3ؾ���(IL����|L�񆺬���FBmj���1�[���@�\���0L��DU���fYq3G�qf�WmA�$����q��l�e�о�	/ötm<	�<��e�'S3����3~��l8��uq
S�p�KΏg�Cu _�v'�زN�I��l����^20�׉��y�Ju����c��/�@��1��k��6��i��	ii��C���g��^ X���r�Vbʴ�^ �G�p	Y�0�����yν��tq������V*��l_{���t�68����e�g�Y�1DVb�c�k.7��.��y*]}��a��y�O����(����8�6�/K͕Y1\62�J�ЌSW���Y]�/����Pu��8���]��m�~m�"�O�Q�����-��!ԅ|�7Y/F�U�޼<�)r��+*ŋM�L�t�K1����m���A�z�?9(��'�4���x�W�rD��+�G���Jd�4�Q%�GS+aVbu/��7�u7���sݒ�%�ĉT���N:^�]�l�Ur�B\�\u�v	��>���](��s2�$� �)�0ܭ?ms���g���"��Y+��llYb���|��b#��$ۆKa�6�H��n�e%����X���.W?�.D��lɇ�w���K�a����*��%	���V�L���;�YśX�$dn,>�6�:���N��]�l�<X��ڙ�uvKO�f�.��`�2ӷ�%��\�>����L1;���iԪp���ǝ*i�:6���>C�4$@�FAQ��x�C��_��oм���
\�{nCI!�0m�������CNzu�d�B�
P(Ǝ����Ӥ?޴k\z��9,�!2f[�\���А��C*�D��8�ҷ=�O{:nَ�n>�r�4X�PF1�~���U�֟H����ܑ��������IA@�/zt
��"���&�j�L����S5#y�{.#+�o�\�������dH(��?X��
aAD�S�b��݁�av���B��g^I�|iw�� ����$r�G���hg�M���ƍ͋&.�V�N�x�;j�gH�_$T��b��rĪ�c�cKlؤ.�C����ܻЙs����-�@��4��T��M��1e3c�b��#��b�Cƪ�首8�E{���rh�9zL�c�ξ�[�>�C0��lȁ^TZ�6�d��y7]B�p1�=BQ��w��9y�N�V���3�㩬U�-̈́�>�0�>�nC�H���_)��#U�(�����Wֺ�p������p(���y��Q<)kO�����F��&�T��Xb�aTB(����6�d�M��c�6vk�03�ۨ�s�������o���q��u�����:�&W.rm�F�ǆPF�T�r��o7�w��xuK��.4ڨI���VG 7�$)��*b���<����^��C�� ��5J�N�ުp���vQ$9�3��{0��a���9��1ҹQ������(��X<����%��k{���=T�,�EHH��v	�bW�[L�<NԬ���7����f�t�������dSEǓ�N�bō���6�>�v���c�~��;ͷ���f̹Uv�"A�a2ۦ�1�q�#����8�:П�w���.�UH�=u��c���z��|�)�R�v�2�"���Qh��ϫu���ۨ7�y��i5��el�[u٬�nm�э	2��N;}�(�`�~�����`r�|Ά���Zf�U4���d� �'7����h�7��fa8e��s�*:|"��"�
n����4xo�y&p��e
��&y�p:�5�?E�	�8`����e�ﳣ'`Nō ���bG�-��2� �}��뭮%;7����i[�,�}�tP���3�]f�n��ɥ�����a���>�k�� `s&3<�]w�锆����(k�~�"tx�R�v�4C�ͯ9a��v6��rR5���/:��>��iQ-��<�X%��`"ڐ��N]p�	n"�YWlyē]\eAYKN��Q��4J���|_�����T��7O8�����{Q��D��N=u���M
�����Jŀ�� ��B}��h��CEQ�bib�{��D�R��]�ca)v演.ې3	�dd+�rM�Uj A�
\1����T���M�f�c<�8�ŏ?�4��x,v�P4��F�����h�I��zP�܌����)�N��k%̒F�U�KѾ�]�ׁb�~]rr-����p��E�7mt%'��$���U�����ƹ�p%
"[K���j�0�O˩JAH�C�S
_�erS�Z2!��Р��L���s�v����w���@�x�!	<ukW�hТ%@�.T8�PPg�g���N7�۝u��.q�Lt�q΄LZ����o����1�]��E���%��kV�.�T2;d5L-^����0>����к�K��Q_X )�#���b&�3��Dey�Ux�ǝv��{[?^/��R�)�}�-S���h�U�8G�B�B�˽��AG h{�T �����y	 ��mI&�7��:a �GpW<��E$2;�>�b}EpN`�U8ؕ����(�_��+Φ`��rp�]e-ѳA�N_�]�KX�]H1q��z��\��xQ��6V�@��xIΝ��i'��ٹ��;<3, T
Nӝ�O嬟Z�D����ֹX�*�L��E�p���>���)�[����k��QX#fMm'��T��d���~/!��[����.fIZ����O0m�c�X�����j����&~k��$�k{����=膆n4!�<�t��"��/���V�G�~D�3*$�k�����������L�m.�Y��*KZ��-}�����<�	��U!6��o��;֊��8�TCV���/p1��5]��2�
8Q%�I����X�g�_�X��,��5���Z+\�~�����g���q5�ZD�$�.���v��y� �5�N�J��w��Y�1viE�7cw2+��}ִF�x`��@	���<_+T���,��T�<��������ϊN�̭6��"g��zJ;��� ՞bZL��sv@�(GA�v%�Y��ok�v�xnf��{�]�<6�!���v�v����������ܴ��G��]b0R �����x	����lV0����`�l���Ghk	��e����AX�tCN��Ʋu@�˿��`U�ߏ���dO�Z6���$��i����`;�z�-Q*�,��k��ʌ�(���-bZ�8߉�M���Yrtw����Gr����쀰98��T���..]9��^{�FQ��un=�Ɨ]hn�f�0LBp�h�		�<�}�J)2�� ��#R%� �x���[h�U%_$8��	wu�Þe��VO���X�@��&]�=S�9bS=�&���6�C��P�����b���U��S��՞܂)��+i�������[6Ù��Q@nS�&��=�1Dou��
��uk�ٷ��@��LB8`����vx�|ќ$�R@5�U����Ֆk"�=y���|��V�^ap��5
{�[�x㩕]��<�@8�;��s�7��������&�е��F�~
ѐ�6�"�5T����׷�	_�ml�^�`y��1Rߏ�V����@a�j��m"lCDC�2`� dT��Ga�[:��<�A�s_�_��Xw�g���~�&I7���Ni[�N�x�>`�Y���P|�	��ܹ��5Uz��֧���%�ye;4m[��
D����u��0�iFN<(�:8V��]�8d�7[���o�õ^��,�Ę��ϥ��a(�
5>��o4A�{�笯�k�V~zn&��)\�{[`��:���IV���,t,�����%Q
;s1��;q�X�/��鼴W$��2Y|e��y?���
�)";7��j-y,%Gۥ�=#ϫ.(���h=������h�9��4�OV��a��]ރ�5e��TX���{����R�W!+�w�82�P�J��D+�u���G)~���Xkl
��(�������<.��41��3,���!�Uˉ;eߋ�e�8�SҝH��W~�X����`o(��N�O
�uG��3�w�MM���t]s��7�S�� 霷j�ܯɄ4��?ݝ�\��|��s�79��$����GŔ}�R�t��� _P�+W(��j��|X �䕘�Cj����z2�gY�}�l�yރ"�NEW
�k�:̴�{s�2r��&�26���S'y?
~�у��Hָ�w���ܑcl��0xp ���]�[*m��>�'A݌�N�/,�c�b��c��h�*]���� i-�41�[�Q/3υ;-&_L���"Ebڒѓ�|�q����s海�Ʈ�L��ۿq�Ts�E��ԝ��sw���5��_�&]*v�t���x��hK�B�� ~��L�Ę�U��$�ޔ����{j�@�����U㗢��~�qRPJh�B'�w6���2�|�_���[��j������miJ�Z����m�n�{�h������j�%"늪_���-Ǝ���@����|J��WuM�I����[�AT���q��n}��Tu�9�(�W�ZNz�:$:쎳ϊn
�WP\?k�1ĐQ�r��vsP��+���!FO���W�����������$T����~w�8�D5�TJ-�|B��Ē3�Ŷ�E�|�{�и�ݺ�}Q�=��-_fu�Kp��{�)�Q���3 �ϔ�($��]�P{��ND���F�"y9z�*�v]"�}�Q��g!u�et��N�*Q�#��p�)�|Z��o��W�<%�T���f�V�����|\/��ii3����א�;�|;P�}j,���1Ff4v���� �U���F/�����v��̴���k2��T��W��I<�α�"��Az>h^A��~*���ۻ��+m��#�On\�֦)� g�'xv�:�{9�d����zmw) о���'�"���A�u#g��f�\E��Gɹk�O�ŧ�b����S����*���D^w�[�4�Uu{�q���V��ӅI�X���`�����b�`�Ē@QB�>Y��
"�nYW���m��?��t��8���P��O3�yņlSE�F"Mm�~�q�k��Mq��^T
�������_af�I������ܐc|}y��͐�b���O�� V��E�P@k�^YDG�9+p։u�t��:{�F�_�B��� Y��k�2N�r��r�&���!%�.��j�^݃�ƶ�:~�ғ)�C�?%@�r��b)Rv[�"Z���v�|[�^pf�	�������,��-ʋ������5[�� ����b5�ϣ��3'�u�|�e�Vi��s�O�.���[_Е0AƇ�;������;�@����p#�f��+Ӡ=V��W��f�`�sf^�v�_ݬ��I�s�mZW�"b�|~k'Q�i�-[Aw��R��F�YȢ;Q��*<�e�D������D����O�@1��F��3��+�.�RY;[��j��K=A����7�����b%m.}���2�|�w���/B%����!�z��pJƞ�*�x4z�Y�'P/��O�&V6��Lg=�Cu�7�z���74�I:p��[g�l�ǫ�� ��e�����HeR\�I���GcI�C�l��u{I��Q;G� �ޭ�ֽ�E,G��I�!�$T���o���ԗ���h�����/,[u�o:*�!����s�\����fb�Z�@�A�65�7����W� �8��6dg�@g�����?`����)�7�
כ%��A6ܻӕ���j�jn�+���ST&�M��>������+m;����g����Σ�q���gɰ�^��&��&)�w�r���lD���ّ@�����±lwD�d�]�Zǥ����� j;/(o��о`2��\��ԇ'�^{�S�5�ޕ��x�nɖ8n)ȝ
e�]�+����6(�����H�YZ�ئd���f����k�H�\o*=�x�	��&����jbVe���CPQ�Au�k�6�b�d]�G���T��~��4�:��3S0�VI������ �[7-�rR�ϥ��L�	��9�t�8I����e��K��sه��?�*٢��t�e���ʽ��C�i�[f]t�|"N1���t�m�r�#�L��� �W� 6� 2�Q��/�g�(�V'hÈ��cէ��~O�+��9׮�1f�c(�����K�o�y���;uk�4�[�J8o�E!�X ����� ����9�W�㝈Te��/i��C�z��36g\;�#g,D�Ej�Hh5=��PmlȌ�6xA�1���a���n�S�v�ئ�g������W�O���u�<u��}_�Ɓ)�[7F>Q�*u¿��{o�D�5�k�ʛ�a�u��=<�f�x�[��������������,�(`�4�_���.��jK�U!P&�}V&�µ/t���~�����o.M �l�-�T�ܶx���;�8�o4*ϰ�/�~'}���j횿0����ǻ��V7���1�Βܕ���d�p<0 �{o �:��;3�ï���U��"eӊi8��o~M���H^��3ԁ���u��'o�%��&�B�	UHxy�Q�AH}��WD��~i�*]=xaA�{���f��l=��f$.0}[-�CBT���^��k0�8:�S ^;���I,v�X8���aKS�/�%9O�Hpe@P:�����(@POZx�p�؛p�Q������B�w���X��E����/I���tH�/]���y �D>���=� �HZ��ĭ0I`W���������ou��-���"��y*Lx3$�	 ]瘿Z'[�{�K���N�ײ��/1n�C�n����ň2N��2&9�$��L�[UDV�kS�}]ʚ82u�g<Tl�J�V�o�_��'�����d�����$:5��I<na�'�M�����9�XC�љ_�N�/iغ�,#!x$������3wZP;V׺����b°@==�Y�������'�|>��$P�7I<����;�t��٧U;w�SL��)�	\��T.��E�On����P�å�+-��8�q'P�3>ZhPb�=�Aͭ�6��Z䡦�E0ѵ��D��߭Ep��͊\E�Hž�e���@+ ܮ:c�&�\0�D����a�"o��:u@ڽF��w�S���O��E�/o2J-Å/,�G��B9Rb� �]�se������d�:��e����M^<_H]7��>��VFj�r.8뭺�$	u�ъ`�(f�5�S�����,C�<PYPK�߃8N,�߼��S�(�mKIK��<�r�;�&��ɎS��=?|����(��y�o�kq�v6q����!$S�rei��fH��?���7�K�g���Ԩ�5�N��u���]}�|�.�%��E�?:秥�ܵ�����z�^�d�*P�X��qa�w���/����z?��mÞ�l%�5<�{���s������c�$�{������E��(��~����[��f���_{ş���ՙ.�!��F�����{��_��ғV��Q'Yf��H��v�T! �:q��V�"Xx��-��,�Q����������v^.�Z؃���Kc�89�
`�@�H���D�J�c��������y�2���]q>��m����_�f|�����2N(���@�Qw��W�Lij���R&[�z�1�~�$'�6x���{��Y�9d�3O.[��ض�M���Cx4D��F����g�k�4+ǽ�60�	���V�;����*�1t���j����L��;�җ��~�O�zK�⯒��<���.;�a]��N�l֐������l����.�#���N�����[n��eW�@�qhIz������{��/F�p������$���� �pߎz#���:W����w�G0P[~V�S��\7xK����m���P�6#�N��R���T����z�Z��K��R7��C�IL��<8+�l
��lX�oT ���n�ܥ��������@�vI���ԗ����g���k?���m�ᰶc����r �����\p���kO�W�L'��fk�CW�AM�ǟBE#O-��Rd }���52. g���v�zRQ�;=F*O��-<m��¾��5�={�c��X�Œ����^ăT,ν��k��?Jfy�2bF5�޺>Hf�e��Y=ܛ }��5ZU�k����2C�Rб>V�8O�}c�?�v7�,|z.�8Y�/|v���X���s}��y@_;�.pP�Hg�o|���S�pk}�]O�����^���dt����}t��hq]�O d��kSE^�)\0nd^�5��̡��,?X���g��DE `��3��yt�$â5�~$R����Vx��HP����)����K�diE�]�:��(���1�����u�J;a�,�GQn���).�({X����r�t4_��®�/��Im/�;����!�?��%�f�� ��/b�c�|+B�r�gow����O���F�f�Z4��_�l��m�?V^0;[UT���i?�=��g+�0se�����.Z��b�U�;��6�Zλ�!�4"[0�g�f�i_�� i6:����ڨ��o��F�%���^�Y_�n��g3٨���8��×�0U�h�
m�D�x��q
���&��7���R�=<���G�^�մ�GgRnt���g��Ʃ|?~��� dIܷLв������Gr�]�
$J��:F�k�j��NL��Ȁk��J�}{�O�.�21Hm�"`i#��N�ԗ������d��*%�.wBP� u��9�ۙ�������-�,���RL=�>���x;G�k�w�]��1���59ꢟ]�s���K# #�Uó�h�[���w�_k}s�i�Z�V�=F�s�t&�b�SEj��$�A������q����F
A�}�2���u6%Y��	��������~���o`�x�z�x�>1F�����'���rS��78 ��2��1j��^}�jXK˅V'�q�O�[�����417Ȩ4����Φ�gZqN�z=6�F�s�$���ۈ?�L�s;��;D�8ĒN��KLY^��W +����GAj��sV<�۰��Z0�Fa=>.��6v"/��������
�S�dCA�W>���@q��r�F%�+���c�t�T�����^���1A��U�gS�
{
�j��\ӰB��bo8�^�N!��UL1���b �45�~�\��8L�)wB�k���m{� �:���CzJ�U�U̢X3Z�D��)2`w�(��H}��kT���O��㓕6�>��Xv��J�B3�`�NN<�)�W�&�7�{L{0�A��AQ�.p�/��+�S�t��>x�Dp7����UJ����Y��SN�jƼ�nlή1���x����d��;u
ުH���֬�m�fST����b�\�U��.���s��tK�ilH����ϐX�\�in25b�>&O��m�T��c����u�6��$�S��9�$t�A�9��ٍthyɌ,_{O�U�R����&���q�j1�U��p��FE
��ƅ�� �����}�4[x;���"t��[��pmmM�5P��v���Q��6d �]�ʚ�-��25j��yIK�΅n��>���z��w�~{�r��i8�-<��~�S����GF�,W�=p�`�~�L�rI�o��78GI@jo�̉��c�9����7��[#\mt̻�i/����޵SE�~e���{��̗G�M�3�Ξ�P�~g�ee��F�n�kA�OL�Έ�v��l#o��������E�<	1���_���@�@bl���#rڻ����rxy�{�e��߁#/G��2^>f���.�;�b�R����#9�Ԡ�ǧQPw�y���z!���mHa+�vvf�(@������ߝ'�n�=@��V��\b�m��㜢��q"f��FfÛ�����}v
�K��:�"з�Q�o�X]�p�������<���>h�����l�$n��;���S!}*���8y�x����j;#c�_��R	�m���v��R1�1@��$��`��%��Y�G��w�y��V�ޑ4xA ,+5 ��������՝�nIP��ф=!���Epw�̲�=s�$�xl~a������4�٢��۬ �f�n��Mp����s�->��n>�gؓ�I�4�?�4��Ӽ$!���v�5��g�	ٗ��_'�jGl,���z����Ւ��^H���nc:��q
ӳG�,��AU,Xw��i����ҕ
�����Z���q�O���o��ꀋ'窕R
mM��H�O���w�tZ6���A~�5����%Ѳ�f	w��`��6]�q�T�.K.���"#�+�8�+����Wpn�R?9r��`� ��b?��C��[�'c���b��SEf��ꍧ!W�i����W���x�?䢆$v+t�Y��G$k6O�! tK���ϯ��C�+V'�[Z1]ԅ���|���+Ho߮r�Op���jճ�Oޝ��˃7�?��gG @�t�Y܊��R��@D7b"��>Ds�X'�O��g4��u���WTQ9C���b_����a�t"����Y*������Qԙ��7��bb;��Os̢_���A�Z����"�EJʽ{��@b@�w��i�2�� a~�1/�Υ�x��,��KB���NA]-�ߑ��i��m��--|�EA{�vwJ�|�w��\��wa�@��we4��=" �[MJhM��U�c(LA�܋2����*�x�Tׄ�΢�d��ۻ^���n�p\��2I��� sg��n`TH9<�p]��)��6���_�u��Yo�s�Kr�jÃb�&�ڃ��Yyב��^��v_�.hʣ�E�mVY�>o�p������!a����Uf�^z���Z��˸깱[�R��]V>E���}�=<����`pc�@n�G��Jm�0S�b
j|��at��m����&��!c��W�DF�e�M��~����r���Y��b���g�%-�_�
�%��+|�ڶu�D� p��d�)�zgL��	X�V� �һC�g�����d!���i�_	g��ּ�l=��)�^3�$�*�ТX=Y�5\��� �����N[E�z�|&��L
v^|���u�?h�|�]@''�?m�bߡ�p���[��u�˂�=x� �f{l�������؟`h'@��}5�Z��ߝ2L�f�	bvA����&�ݢڍV}�5I��Dz����"W2�%�,�>݃���ۼ!�-sr/�*#������>�9�S���q����n�
�~��6hW�������}���*58K]��Y��뮞��] ����	�O�Q�+��������K��.n��&*�M즠��0՜QS��̆�TL���s���l��-�u5?���|��x ��U��w�	^}x1����O4���*�3�V9�1���zXr�P�A����ab�rwIX� w9q�O}���'Ҿ��m�EX~Zu:���S��3�k����������ّ����]Ҍa4U�D9�JP3\UhB(���xo��PpS*��4u!Z�ͬ��:�(1�gI�ay�`[@!�z7��n�ª0�^��j���v�Z��A��>~^���= o��C5�wy��<)��i2��wY]gڷ�Tsv�B>z���1���Dg���h����LL�� ���|��j/S�S�-d���4>��坑��+u]�͹�k>.Բ�y�P&�j7k�p{�\LZ�zf��ej{�c��Xk�J�%���-��&�J�%�[!������N������M���{^2`���o+g�f�x5�>�7�/=��)����m�t��%0tg�^[��;�Z��*�`�L*A�Z���`����C��q�u53�NXذMB�q������~�l�\p����2dQ:+>c_��L���_�_�u�b�<+�<j��A�%Y��1������R�H13k�^��c���9)�}�Xw�h׃\Q������M�D��Wpx�5��~��g��~"�v{x,N�6k`��z0r6u�b:�K�š�(�9�jꂇ]H��_����5�~�.�B�艡�y$�T�y�o,����~���v���2Ҙ7O��Nzy�wi�"g)G�/�V�صpv̨{�f�N{�2y
�jc����!GA�4f�^���ӗ��}'�K�#aOF8�[�L�{p�^/��k���{�91� 
j��K'���2B���9'�@JI�����[�[�KV�������%��o��L �����ߋ�f�w���\eg6�Fxw?������h��{�$9���Q�4���1�PoRJ����g򹏆�ɳ�H���eFӴ��p�	�ֳ���:9�x�		a/{����Yޘ�i眂|f쒈��� pE.��J�̞��1i�v�Ot��ng#�����ë�����Ѧ��,��G��c�-��Gic�+2����~��U�Q�Os��Ӱ[E����xշj�
ʙW����yoz�H�_�h�>�
�}���L�����ܻ��H�5`��DdZ�#���7 �W��F�=g���X��cT&a��=S�0-��o	�@�}ӱ��gb�n3os0�9W�eJ��b�V-`���Ȯ.�uǮ��qK�|��g��B�}�+�ч3������q����` �*�C�p&w#�����.��
�y#��w\��"��F�y����� k����̫��(h3ؼ�P����d=�p,��~�qB��9*S[rS��6x�{{�о����j��e?�)�'����O�B��O�m
�0e����M*��sW����]�4��E�2���(=�ݺ�&iq�5���P~8���^#�Oy1l��1��C�d
���t�Md`��b��c�h�]<���v��F��Α�V���$�
��m���#7��C��Q��Ύ�?�Rd�3z_��,gWre�Mk���U.��Q�bC������W�.�G�ڋ��ю��U^�e�\�sM�52�.��o���S�؊�Z)��~�T0�e����7���[�&*[po,�EwD��p��Ý�ߓ������I��;nB�ҿ�v)�C*3�Hvaӿ�wS�'C�i�)��Uĭ�i�|��;_�C0N���Ƕ�$:.�P1~gw����S7�H�=�3L���S���k�Z;QU�q��s��LH�˽cvoԽ������R�2�Ue����]�u��L�?-�8�CY���ʩ����W/�U��þH��J�>�~1b�ވ����?V�@M���?��e��Ȃ6�&��$�]M�/��&%���у�eD���x�ٍ�,a�pݳ��oi��?
Y&���g��7':|#s<���]񜬁��׃;��ߎ{@&�	��?0<�}@eBҺ�QM%S=�Qz���%][0�x�i5���?�\���0C%�_j�9�&�(.�8���z���4�]�O0	x����ٔ���2��L�����K��ɐ:Kc�����q�� ���SR4�m:�_^���~��)��߿�9-+:X�ά_>�����&>Y�jR5��b�^��m�EL�+����y�� ���j�W ��^!g%�m��+�y���� T
a�Hͩ�����1�մl5o�������G^�w��A�<p5�tjl8�۴�aLa�)3z<'�v�W�����`aH�Mc4�t�r�?��R��ʶ�p�Ϋ8Pt����3��H��V��z�3�I¾i�+6�pG��BJ5Bf�C䈢�`�.^[�����ZE��ð9����pZ�/���QP.����G~��S���9AQ� �=y�cwF\�����4	`9���
��Wy�
���!r�Y�3 ���ݎm_}2T��ia2�==�7O��u+�^)F X����x�	߬O��p����ٛѓ��.Lh&�I�s:�S���ߣY9N���4�<a���Mm���u��hiF�:MAm b�@?v���ʹ!���i�\�x?޵�Z)3o���!�=*}��u�:������3z�E_���[N���đ}At�����%Ӗ[�Jo���ã�G�XE �Ȣ�	&X��o�Φ5�����+i���ӟ��fʭ����')�aJr�=���=�+��fgލ?Wa/���*�k+�^��α���^W������ߌ3�G����E��T�Y�.�3׌n?�ϖ_��l�����Z��8-���[���{��x�����/P��bx�<9R�b�@D�Vh�<����9� "nv��3qvu�ׯ�=9sZ_ .JqZ5��!ipȳp$�¿չ��b���*����/���s�8�<������M���q��RW;��@�����Q�c@쌒��r͛�p�k|T��7,vo"I����U��(q��qR��WJ��ܓ�':` Y�8;��b�2��vm[�tz�L��]����U��n����ڤ0U���>�[��Y2�⡦5�t�~��e�$�F��UJ�={���������'XS~�z�ȟ_ȡ��۫1~'����?�|���(��������eT��s��Z5�0_���t��ɇ)�ݑ�px͜� �pW�Ϙ��\^��WuG�>��t�O86Glƨ���S~C�/��3{\%�aw>�VK?O;5P�[F,�@�SCc^���ta��ǖi>��T���Z�����w��v��2+�%b2��t�=6�	 �sBpw���e._>;�qf��M}���ch�n2��� ���-��͡(Q^G��C4�{� ����&�d�~��8���x"�7��z�#`\�(�G��a2��R������!X�/�u�`V���G�8�f�v�Jt�2t2>���e��ƭ#5�&��Vc6l(&�M�T[�~s�z��}z��
v�vk��� xAak�͌��a�:�OC�� ΄�]�Czb}C��뀻π#��ۼ�R���~*_YOx���Μ��FXj���=n�?+��d~����<���4gO���E�l˂����Wy3�I7��-�(��Z�����	�=�$�Ļ�P�}��o��^�PJ�}(�"�V3=��.zh_u�P�(f*������"�.��v�p����L��7d����ywė�����{\����]���~N���z9����������Pr�y�֕ �?z�ŀ߹Ǘ%� ���`��ǀ� �	���_�*5�u&t��G���7�ky~�5�`�s�b�#} �`����ꥺ���c4�����Z�~�T%��$$�˪IM+�)�I�^w���?3'~���f �Rq	{�c���B=��Y^��;���X�Y<ʢ��F�� �b�Q�40�������
C��X깑�>�� �9�����f�g��:N���M���o`�  ��Ǔ��-�dN�b��j.�l�{�$9q��L�� ��_��Yؖq`�I���lC�
��]����$ዡ�_�:'�����O�4��I��q�g�b-���F�pOv/'�yp��?�4c������]]���,_99^�Ä�]����	��MQY���:{n�IX�9���p��y�Ln5��i��M�4pbI8)|7���;�3��m��7®�^����3o��9���a��l���u]���IA��t���NFܸ�b㥌\���;�4���I�6�������+s����gO�πr��EΩ�Ky������������f �$�u�/`�UN{��\EH�|c�(���^��J�s�QqB���<�!�XyWpu�9.��O�`1��m%�Z|�T���tY�%I���e�����)q��6�e_յ�IҰ����-��w"�bV�&b�Huy��/��'n�ʥ��ğ�r`1|;���)��g9H�����UBp&#�-�\�&��8&7��)�t���n�^Rs�R�#�<K3���ڪR����x2������9Q��]C�9�cܣ��H����o�YQ��o��tH��K�Z����b\�r�ҿ[n5�ۂ�?dyaΎDT�9���/�ڿ�ɽ
*�#2��u�
X�?A���c���x���������{���(g	O��j����c�L�ك��܅�2�$��
����by���<g�2�H�H��㉲nI�����,BЉa�o��rA��s{�4��ѫÁΩ��c�o��@����ޘ;���#-}�qP�v�D�!�8r�f2U��wH)�鎮�_�ˀ�1�v��U���^�q�%%���?tȩdM��!s��Y�p������Ux��ܵEz�����_�����#�[��y���l.��e���rS����n����f�ȟe��������eg�#�̛�D����u8$�{���d_�.�ۜ?�+)��)��s9$���"�6����?�$v;�۳����ɶs�����{��!:@���I�j��@!żc$R�}�En\
Z*�O\�y�b[[os�u�Q��H��;�bC�А�Tk$!=�GOx��Q&]��I�0w����vH.���n��s�E�&�2��h)�����R<��c��0������='X�o�4#�{�`%б���5V,j�r(��zZ��ј�믷<��%�¼���/i���6���W�u.�Q���?�q��$�lE��"va�_�
������8����M*�/�Ҹ�ZS��*J��BU<FIw�4&_���?y�G�αS�n��I=}�
4q�ʍ��{�v��c����QMvx."���Z���"��L��aȍ2["-b5��:	�c�	ۊ�?uH^�N=W&۱�7I���+���=�W�c���*�ׯ�6���Ȃ2�+��P�����K%j��8
�������ɭ����ݩ����:�la���*||Mt���r���.��

:��q���ԉOBG� %�K� ��G2!_���<��p>\`S7U1X�O�>�d�T�|�t� d�s~��������4�p�L'�����NxY}��vt{��D�l��l��>���,ݛ��{4@�o�tk����~^Y%LHf�ࣇ>v?��Dfn�qÄ.4�W����k�� ���S{b����}d����p�߰�s�6c�"���iZj��A�k�@Ѫ�����A�f̆�Mf�>Ҍ&Ӎ���7fX��C,�Ml�o@��	˥���՞SK�6��gT�E-�Dk"��$,��a~���&E�Io/R�{?,�.bչ�!���uipuԨ2�Z{qs��˽������t?.��QW�^����~��mDR�_#��Q�\��(�����L�7�ٍ�߹��l�=H�ş����q?��\��9x�TjX��Kk5x�ZM�e����KL<����Qg�zW�G5X(� ��1�U-3�+Q�n�'�$�O��h��nB�d��k���Z���g.���	�����.Oo��,��54��[x@����@�tJ��+�����Uj'�G���Y{�)��׍�q��Z����%1Q��ܵ�$KԠ�s3���)�4ps7pO�m�k�i�te��V�{��n���i�w�����X:��T�&WQ��FT�:����#�}va>՘c��9J�ۣ���4�؇F��MR�v�Q/'��u����<�� 1�>*��Z��u�ݵb-��Mg���H�P�U����1�1qR�� j���m�iA؉T0�E�L��_�,P�ncCBO��\���{�"�of2o�����j��j��w&�y�I�@�ҩ����;m��{ޣk���R�2k0�+�d�|���t�(���;) ��E �/���@�-@�`E�����u��l
z�"��0��ܜ���wu.�����K��w���Ϗ�6%�P����Һ�J�@��Oa�/���d�6����n�J�'�h�Y�XE.�'����kJk.��c�<	���ys����^����Fi�t�U�&�+8�.���pbK?�1| Pp��Ϸ����!|���ɡy��iCBל۩7���7���\z��G]�d?�od�b�ht�w��\Uy��YR�׏;A��^�(ܧأ
����˷�:׮����u`�,ߒX22UY<��g��u���;�+�Յ������3`��Qک��턝5�>;r���~�@'vx�0���^-�W�W���~�J��`_�=ޚ��Vb����7���P<%�2d�vq��J�D��{��lT��l8}?�>��.�li�1�q�yōVk&�/=����SC
�㫋�Akk�/��{
�4��,�I��!�t*���0[�n�� �ϙ!���D�.M���� 2��w��F~�^v� �n,�Z�Wh�Tc9����Ro���+�!kc����,:f��u����#����-|p)h6�/wY��ud��m��J��V{��F��EӨc�t��2AR��\$.;o���T�thӰO��~��PK��ҥ�-��ҥw��
~�[��?0��M�Y�+=�;�U���B��MW��u	A@��.�RA)顑i����[j$�a@Z�nA��$��c�7��K�b-]��{�>{�sߛ5��(ѥW��	�Չ������n>�T�}�`�wg�?�v��'G��J��4�c+k=�BUa�˓�/TP�2�T!�� \���fY!��;�P����}!�(�?��_�Pn�1�����d~�OF�08zu��YQ�	*��P�p�߾ �>		�%�"�������ػ�N�18h�.2R!��C��o$�����sL�J�߁������7�v��w�'� �ޫ�Ϩ��;����m�=Z�[�F�.\�1ᡰW}ZZrw��� -Ş�����*�|���]�S�J���Ki`]|�6zR�ʻ���v�NeK��x�}�᧿��NZ����M����34���-�Q�h,�S�����-�����s�Aˌ�J�jɗ�L��q���c���~�֑�
��T�V�����~N'��O���U�g��d�0�"�8��#l�����c��,5�M���>������id�Czϭ�Yr׺9aZ����s尰TM~�kc��}(�$��F~���4�rf�l8�1�
�r�Ae��O���ᯰ�*�󲯻�ǚ0�.}��:������^M�/�㵶�����!��KZ?����7���&~l�ՙ��u����dH��Lf��5j?�RP������=�j������7��
՛�3�q)���6�V�2���7�]�
�,�tj߄�M8*m�Mj~�QW/j��(�wT�ؙ�,���wPR�@H)(=�o"0���S2�N��o�h�ڂ玏&Ֆ'U��hY�5P~K��%|�9��<�w�J�V�����D����_��8�C��:����}�[���*� �������W-l�Ԗ���HB�K�$��~&� s�*b� �P@��v]u
�=�	����R0�����I�׈��h�_�֋3n�3jY���G%�E+�}κ˒��jE����X�Ǘ~�ϵH�6U�4i��\%�������T��{��=����K�-�uY�:��9��y{U�J)��2�*=c�u�y�1�}��1qk�i��"�/x��&��y+������o��V�����'��}��q�cm��9����c��'	y��6�H�������f��m�8���x����qx������şks�c�%���Ao9���C��*WyD޻:#_�~m�b����Z$�C����%C���ܼ���X��?�5K'	��)�h�TN�p�˱@��8�~�hp[�dk��ӎ �\����-��ԤdZ'�r:��1̭w��ӄ��xA���"FTg��`�Ga��cO&��E ���1�t(�j	*�Q��V=(��~�F��c��_WY��ȥEGo�Ɔ�����0����4����}[D1"��+�M�T�=!�Ԥ��=X�BA��G4� �Eq5�!7�p=5X��[z�`<�H���]��$�r-�zC+$�6�)�ͅx�����-�.�t��9��G�*;���&����iO��:u�3��!��o�&z.N(p^�d�t���?;�P�4��s�N,�o(�#)�u<y!8���2b���܎8U���a����aW� x͹����4�p)u�k>�{X����t�l��,��h����13�YwQ��� uT�� �֟ʧM�9����$uQ^���M����|��~7%o<c���\�2��,������� �4��#����-��ţ�]�p�7Ob9'��Z�O��6�0
U0�'�ʙ���j�{�%��8���F ��v\"g��/U^�y]t�A.�(OUQ"XU��, �nq�ʛ ��4W�(3z�psM7|�̠Q��9��Aj7S��'��`rxti��uzt��DF\�ު��'n���ݍ�"}�s�⎁GY�u���~�3���¹���}����Z�8{�>��\�_�	Q�������)mz^7i/ z�ooB�#}�ɇc=�́<{�:y$2�뇳��,��/�k����F�b�IK��_ٚ����Y
�hq^�?�� ����;�'����fug�Mm�.�p9�*C�4�Og�/EW�(���#O.�
��:H��H7gs��j}���j"�\q���������
��8��JT/�FYpi���x��N��	5��ݔz��̕v|�ﲱ>��n�[��r4�ME�vq}��IȦpۦ����b\U� ?ya:���f��ח<�Ҋ���[N@+��$�R�Í��|�03���O��?�Xu LN�NYf�Ж�����q��;�f]��h�h7�%5c����r������i���;i��{�N���8M�t��/"�Z}���	���+�*
N�gW��5��*5\�y�oƾa,�"��̋v�>���="#kY��1�����5�u�4�]�&�d �l�]M�]���:��:����d�2v��d���8�?!o
���fi�����V�X[�EWa��N����ڠ�VP����(��S�Un�����	�,��K�G��]���1�q�{��4#zԓ�Q�ĭj��vQ�Gk���)�HO껸\�>�y%eUy��$���&��"�`����\x�KY��S�|f7c���
+��;O��e�n���0�ZĖ�tz��r���*��l��䦝�fl+�,F���X?�%�#���i�s���sS�O�t�y��2j��ʷ�ſL�ѝ�"ܥ猝~j:3cH4�Q1r��h���B��s̠���<���9S��C�:��z7b�t������#NKobF�$s]�
��H�u��Z�$�i�V�z��{Ֆk۴,���_��nk�����ĤM� >+�q�:5]4FVɫuu��x��3d�g�N4��]�*��e��6��'\~dx}q�k�.�Dݰc&�.�`!�Bq9�"nD��+�X�qS5�T 1cN���XI�J��ʗI�����������q�s�叢�-�m5C�Be�"GQ0�L?����Fή>A���R���7��-��~oXp�Mp�\gY��i|V� ~�B���m���4!���2�.=v���_Th�;�߁�;"7Y6��\iBe��Ro�[y����K�x%rH*kJL�7e�|V�rJL�u~nh�/~�,��zGC!�W"�P���������&|�������4ކ�^��8�)�J�ئ������aA�Y�ig7��!�sW>-�$���W�:e�����ʙ(���S�Nec�����)���'�%`Y�u7��Y9W�����������q-X�՞~��x�-a��z�0���R�����4��ۚki�]�dd������7A��k5"9�N}%�9L+��㎷lcPXa6�E:X�jf]�;H�P�	9ŢU,횥���>2�a�X�n�赭�=�K��L̛[ΰ?����O����Mlc�q��>;"㕘n [�M���N�*�l��F��qU�fpgH'(�k�U$l��a.cI�(�C]A�'��:pXYJ��DT��x������uX0��8ׂd���qdZ��������/+t��:�133��}��$��)�
ITC�`̅fS0�/n��L�x��@cM[U�3H)fr����l��Q��7��Kx��� !��T�/'�ߤ�E�R-�H�ȧ��!�]Ud$&�Q�h���s��;�����5#Fvį�<pΑDYQ��5V��W:���A/�Kδ(�|��({��)�F�T�.���l�̳i5�j=���c��QP0�\�t���k:��bY<P
�/\z��M���o�@�5m�1��J�9lKW��9��;W�G�B��ia�_��1�����o���@�G�C�����t�[��I��X 5q��F�ŉ��
y;�8?�L�[��A�>bn<�CD�m�N��6����L.,a��?�F���<3�����»�W�-�t+b��5�p�Y�Agfd�a;�c9���3;��R����Vˎ%"���F�-�һ�Ӣ��	��Z�����l���Uc� Uɶ���b���xx�!p9��٣�mV��E ��#^�\z��	����VK=���&gǃRB��k�Әc�J��|�|y�_��fu`��vT�|������$�rr���d9f	��˷�h��nn=}��SQ��{�M��lc8d���G�=���;�塮��
�6�T�̧�i#n�3/���5km��#"���i��Y������9�edRz���!�R�˟���6/���!�.�R�1�O�������*X#\��f���6m[�ݬb>	�1�}�z�	��y�[���{6����1���ͭ��M�i�U�c̯l��	[��Z�ү�n�z���z������%|��6��5PP��&K�!7F�B1�Ϝ��b�76_��_�/IϪ����7����,���h��!ϯ�2�?��,佊c��:8�VP!������<�B��;C�K秹���Wu'��c��Y?��?��%���<o���tmsڅe�vCb���/�>/�~^�����&詾����o��9���b'�SK�����ʩd�<unt�j�\�?�˭����u=���0P8�0U��)�������浧��uWO��͜���y�C\.�㑌Dk�l3w3�6��%"]2��-Oau����.�Y�f�A��E/W��������	u�T"���;o{�ay�ݍGų��+1���H��Xy��}������f�0%KJ�;g�Ya��)c���+�k#�~[�S�E�B��4��z�)�C�l����,� eu�G�}j�����e�j����B�X�t��REnpQ�9iXZ
�*���f)T�_3zNtY�"1N}hs�5�����@^�F��PM|k���ʒZ}�}�U��)���{���W%�0�$ҷ��^�tb�ι���{��������"r�e��(��v"c����[�F��1��/h	�/��l>N�>`�\��Zo�8�f�t�n����!sȸ 5itҩ�B䓾w-��(��A�Z��V���OM8R�0�]+��ɿ'�I���ʱ M6��q|q�_'3��G-��ʌU[� ��P��@�Yd�����{���臵��Pl��c��~R(l_"���"5�U��ri�J�����`@\7O��4��S�\c��� r��4ĺk�-�R�;uy����&4[���Qf]m�x�[�dw�ύj�p��{4|��.j�j>���kK���]��Č�7S��~�O_ˏ�I�O�����N�LYI�y�	|i+�Ub��ӿ���~��a&�_'u��������{��V�^�`�Zw�)�Z#\	fQ� ���F���X�s�𙆌���fw��5K���o��e���n��x�]⨅a�ϫݕV܅�h��0>��v�څ�ЅP��̘^O��q���D��^k_��_N�(s׻~�C4�H��;��o�ƍ�h��h��6�3���D�r��Pp�s/�R{!�k%�8���O&�`&�Dӷ��6� 2��s��� ��42��k��A����;g�c=�-`�GF��8���քQI
�8P���jN;~���'^p!�>0"$OF�����)
<��XZ�����H��<��@8U�QzA�m�d�8ޔ8?W�!\�>T������Jx��=�{5���x��P�v��7�=�����oPf+K�@۬�� �,���z�RK�Y�7��k"�jk�u�'�psc�ϺwP��R!��d��!�lŧO�DL�k�&}5ږ�nI���@�$I�8(��*U>��c����xZ���hғW5��t���#��j�_$b�`�ο�;l��y����2���p(��E�5�p��Bvl.U/�h��}��az6�B�d9�3�\�D�^��/T�����G�9�
�j�ނ@P��ަ��g@�x�K�4�!���[	�3�r��IF�ln~6#��v ��?U��;����o ���ι�ԅ��b�%=Pd��,�$t�(�t�`��P����8�s������;�%�
 F˺e�-�K=sU�̦IT��/헲�ݕ� D�	u�������9�SH\��H��#�_��</�ʏF�R�̹;��t��Qu�$}Eߋ�mi������4mz�����a���&�~U�Os*��#�����`/�'-�PT�"�5��
���	��Ŷ�F���%��}�0�?`DùA���Y�͜�����G��?�<Kv����!�@�0ӯ���B�}3Z^]��N�Ǚr��	�Iu2<<��;J`�R3e�Nܑrl�����P�d�/q�OPq&P�-D�V�꙼��'�d�\ ^��I�!��)�g
��N�dAhWI�2�WW���f{k�X �c/�����ן��̓���sǠ<@<I��������ڷP�G�G����O��&P���Z��[��i�5!��h�3�!�>y��`���ꌕ9�w]Y��s�Z����%����us/M�3~����߇�E*渚0+o���3:)Ф�ٯ�I"�(d�tK�9 G�ur����ކ-|v`��IB�"2,��KZ�:��W.���h\D�q�i�&�I6�W��!�ܓ���UQ���n"1sU�!�����BR�������m5oq���P�=���ܯn$��f����9���(�Qr5��"��:�z��=ܤ͒ %�#�41`�|�is���"��bǸ2�e�P�a8��a&%���]J��Ռ��3D�ճ�H��l~V��d�0�i�Q Mr�=ёEwg� R,��ci�<���q�k�W�����Cepw���[��Ӣ�[�L��j��F��"�nG����A��Ůo�Zzj�w�e�E�����7+�g����tF�1�֡ݰڊ�dM����ۢ���3]�_�������r^0�@�\��*���h�t���3=�:��ߐT�&�����ͬ�(V�̰Ra{�5��!��wtCDS~�� ��"S��$�TSǱ�nMa5A��>8$I���_,�uv���chY��,���Y0����-O$g�� Gi�~ǵf�ł��� k
��L�8��6���)4�Ѱ7\U��x�3�Z�C�b�S��9��F�4�8.��ߔ8V[�q^�K����� �Y_t8��Ւ>�j?V�/d4ۀ�{]��U�3�r�U�PÇ�&v^��kaK�oH��6�k|�| ,�a�0��}��>����P��#�F�+�
���X��0�n���X���&z�Z�W���v\�/9��
�|I����~�S���2�9�QFev����+tS�C��6eZ�2�����!�DM�ӏ����8И7 e�d~��{�M��E���%u�w���W�[�����e}8�?���r����l4	��P��m��o�W�f5n"��%� :�-ɗf���R�}�� ����C��}��]ޕԭҒ?��U�_ �Rjy��SZl� ���˫��$�n�L�e:�1X�
|��#ʙ2�Y�r)�g��[�$x^�Fo�P��{�j�`�5X�2r.�����>���0�����ȶf�U{��x���a��7q�s�=�HP��(^JObEi�����lb�:F)��9ɞ��B���:��i�&9n�*d4D]/��E�D��NW�:{� 1�H��!��|�Z��!3��(�d
jA�Y
���`�h�^���}Ճ���cp C�c=�fF���3-��9Di��ɆU���H!���20���x��?�B���Zr{�l̒�&Z��HB��Ih߾-���Fgt{��7��sA��s��	<ud�ʀjٯ��.������,�*�#���g[�*Sa3y2W��<! $к�#����R���9%�큞2��]�m_(Y����6�IZ߼k��ɅK3�҈�/���o��ܨX�##|��8Z���
۾T8W�	����Ң��{�O�\��M}*�Y*|��檻O"@�9+ʯM0b�<��]dJ��m�%Pf�ؖR�l��un
lO�<��bN�.^6GĘs����F6k��ehv�Nh�)�0������沠�<��>!�v,@�y�r6k۲W)�XZM3�*�v�4"?7��X18���q�infPjd��7������ .,
�aVl��˺G{$�pb�����<�CML�� �Q�f��o9�ǧ�V�̏�9cL��@x$S3-HH�rqߴ zN�GzI'���\�/=��T뛼:2 a�j��?�s4�`-���nϒٙÇĚ�4Z����mVU��<���*al���$SR���X)z�,s	�^[y$Q�+z<50�#��w�F�ȟ"�_�l�aJ���]i�,��OS�NniG�Tc�~ �in�X	�p��~P9��3���R�"0_��O��#��y�ش�o��ߢ2�?��s'�㭟��L:}&���u:�Q�i��(`��U>�*��m��W��k�K�1?�,��c:X���hD�<7��8V�.��:,��L�N�� }'("�q���a�|M���(��I�mڠ�!ʮ��n��CE|3skp��ds�M�l�!��8��bG��y���L�h��<��x���򼤸	��-�BE��a)�~9Z���q ���+�!�������M'5NJ�#��^�B"����xd5N�*k�aA7�����|^���8�_��"?~#����ml�uE~!ZZ-'�d�B�?������#�e�F�7福g�g���t�R]��A�U̹��� ��wh�pm�;�9\�	=�w�,6
*oy<ُ!�n|���a�cA��|r����?�����g�vf�����"�����S��ʄF���bΨ���2�AO4Waƹ�Ew��1&��q�	^}���$ǚ�`-jy	��%,��b �w��3��1BЂ���NtT�L"s.�s>}��^K�,��U!舰��"�+�����{ph��
�G��9�vc:�˹"~yBw'��+̽8�9P���~5�J�߱�#r
L�]����$���\�T���KLp����D �8�G�x��Ma�V�;Տv�.4�*n�#����r�YW�{�4��՛���Z��X�Ԍ��"�)����FE�"��I��E��K��!M>��h��%f��	F�9%�ܿ����G�>/�E�dH���'�b%VQ�"램������8핲�*CU�u>���qJ�Ez�xE��u� ��Fw�����s�_�>�0��l�\�^���^��\&���)�9�Dͳ��~���3�˟����h�Τ0θ������(�v�X�c4�j�|5�,r���>U�.6n��NhB%���M��<U�{Q�����Tih6��1�E�'\���t�,%@v5&c�����5�:=ڕ�p�ΉT4��C8b�֠�T���_�u成`0�'xy��մ s7�H�LRI\��
�# �m d���G�+�'8CB#������8�����)m�/�1#ၟ8hn�{�=N���v���gX߰�G�/�$'[�%f�}�9LT�W�+$�g��J/�Ev2��mԜլ/.�ZE��C��
5E#�I*��%�'�W��R"_IweT~ ӗK�i�C���7������ƕՖ���p�zT�[��(	]��mϵ[�c�h��%�I��߹�����vQ�bpǏ�]�Խ���t��[��1ItBU�,M���(���Bb�(6���*���c�܁9RmB����`���,�赚�s�l���4_D��G���9c�����G(_��۴�Վy@�l�">���a��*"�|}���H���F
"���o�0FPӷ>̑xRMCjÌL��ůA��M#�Uq�9��%D6ʹ=��{��!�F��.2g?(��2B�������s�lzbTIW99�/(�Wp�~�x6ćņ�D�Ҳ����븢��8��A䧴�:g��\�%�'8u��OczWC7ZC�mw��6?�D��>6���I�iӾ୑@p_Gh�ذ4��W����Ѱ��VDU��x� `��O�����=����o��%�=��}�j�_7V4T�N�NwW����xU�e�/}�:�����6i��'y�2�U���7��
�h6�N(��W����u�8��{t��s+	M-���#�>`�<�d9K����=�
ì#<�(t	<sj!���	ڱ�u���	{ ��r�WU���n�`���D����pP�u]���)�`����C�2}�~�8�J��Ū��+q�pS���ja�i`��v��=�	�~%{w:���~�#��]W�'��ލl�
Hc������M�T��__	+�
���mc�F-)�TPC�`��|����I5=�o���b�������4+�v�t亢M�?4�<q�u'M��U䃳��&�p#����W紉)��Z�a}:�!�8*�Ey2��7�¢9- ���,�����e2����I̞]����8ώ�I��?��S�K֗����E2�~¹��}�Rg�[-c,���k�hj�+�m���m$0/�tF�7�㳫o�@�nU��f(�su�u�cZ����׳������v�b��f��*��RjQ|ÀL��5������v�?��@�A*�k�ȠdE@؋,�ج����0u����<`�s��%�Cm�gU*"4��V�/߈��<�ʭ$:��~���&G��wl�FΈj4�R�q|�\c���|G:��\W@e��;Dz����K��M�gG�a5�]�>ڊ%�8��5�q�]Q��oTl�ohq���u|�RF���A����*UV��[2�Uw����ՙ[����L-J$s.N8��"�N�=�6"s����a`�0�_�sʬvڈ�ctb��
$^��ʗ!�ۢ�GV��~��7F��xi�WB����@�n>1x��WOo,r@o
���Q7({=�OA%ژ7�Z�-��Y�-���t[dR%E�P�����GWX��ٷ���]1�B��G`w��,�7��ߘ������q�	g�0L2�àQ8��	
���\ ��>9nؑ��'rris���c��|GQ�����G�Z���#˾��-�!�u6u�����7�y��@���� in�*��r��Hx�! p@����1�z�!N��n� yr�A츲�B�n�o�M�{���s\U��Nn��T�dͨ�t*���h�p}Ek�~�`dŠԿ������0s�L�ןp��u��@�g!�Oz)�.��b��6��e�R�>���1P3��H���{L2�c-�z�Iq�/@:�-R�DTkbS�z�C>8��|JJ�-mHdwq�>Ρ2����Us�a�>�Յ!���,��wP�+�r��9:�e�dj���p#�z8 p��vr_wF���3�u�u�XbQ�~�rDpE߈�%��4����Ć1�u�����KC ��+"�ɶ��P%R��.�jJ�y�8l���Y`��]��A@"��{���5�q'ь����{���f�['������:��T�^g/�C�?.��Q���>(��������:,m8@��0��u�0dP��S{2{M��Q�d�<S4��iH6"L�
�V����}�ވ�2 ��d<�g�99���gk�i*B2m<QO4 E2���=��������>��4?��k+�S}��
��{��p�j�'����iQ�o#��W��ҡ����v󞏺�s�qI�_]���f��@��ܯ✘����ʸ�܆m(��n�FɼA�v�W��sz�=3��j�{�r�{�ՌE�x����
?��������`�1�I@ �Q���B���{�����Lq2�u$L�4>}n�3r2��m�atݍ#�Z�����M��E>��b�F�Z�mN5E�� F�~���|]��A뱑���,�ܢN�T�?�yH߁r�����_[w����@�Ų[]z����." 423�%Py�
V����픣�Y! L�;�~3e5Q�W��x��"a��]iDq%�����gC�5���%X˨g���`pL���7�F{���o=�{�ĸ!�Ĺ��`c�o��ߤN��Ο���D��l�Bə2�ĸ8!]3�M�a1����S1Nmߗͅy���"�n�3��?�$��:�o�k�!��O�h~�F|���ﴘ���l���ʏbp���/��`��-�E���˟G���7��d�����E	z�7/��!�r@]�����ڞ^�����z`����s��7R��F�
������/D�#��&P�ve�:���0s[$�x�5�?�W{�lJ-(��<H��x�����*�\-r/Qo�]%��0��Xs�w�M�Wx7M
��!���Z�z�9٦�B�{b��3��l�׸��ջ��U�8&������/�p��y�1�R��2Cj���!�"�ͯ���jE�CtxUg�Fj�)�f��JV�U$t���2x���^q�^[UGӻi��8y�9�<�v��N��)�*�ן���?2z?@�ڋ:������M�=���T�՞.H%L�N2�C����������c��,���'��n���>�|p����i*�Q��!M�Ja��s���v�Qץn���a
�g�����Ϲ�=�å~>�"�6�X� �s���~��� ��M4�F�c�f(B�ŧU� i��S���+Mk��K}l�#��[}��dJJ K�.����g3��m.(��7�u��UYh2�����V��(֮`>���)):��U&��ぁ�nW^����D�G���er,�]��u逤�\ kx����.����ᑕ�`BBG��aӻ8��R�g� I�ҺK��z�~ߟD�uuMh�'��n��ɪ�J�p>+�m��E��>��������9��U����5y`⥜�4~
��	�x%�����NU8�����_tW��P0/և�ſ��	�pv���3"��ߑJ�H�8o}[ޜ�ex�`+���|��eyJМ�&t��gl\��kӥp�G��S����z+1�+�%UE�uG�̿�X���sL˅v8�����͇�|M��C��%�}!]��}�~";�͖���5о$B�����*0w���-D��ƇUkP��[_�T�Dn8�Oo��qSȪ�zL/���qe�) �f�
pMzޮ��j���ir��շ[j��r+4�s�ʧ�w�2mu�0�4$O������v��h��n�ӯ����˞S8k�[�J�!!`�V�s��)й[�4X�g����C����W������ܛ(���.�2<m��}L����)�i���0��C((R||jny��2)ng�x樛p5j��&{(a��5o���/*���.��3U���u��U��]�I&��w1��ش�����Ɯ!�\�1��v�E��9�[)��r�K\*%��|ch�zuw�C�#�&��]lp�ƪ��UW������8���lϿ��ӻ�Nmvu�ϧS'���e�0�b��؈���,a�"�MK��R R �3ez��|��B�+)�]�Y�`vXk�_���p*�� !�;Z�=f��;���<_�?Rh�(�12:�@?y�4��7[�d9[�#.3|f$���`DLr@�k|Ԓ��.��zB�5��5��'p�f%
�*�V�}�4���
�_�Z�0�97�u�f�87H�B�e�|21k� �/��~��9�}���M��JVģ����`.�@��ρ�O��Q����X��|�����'��Uk
iL�#���~=�a�n.h�>��( q��꧍��=z�xFf8:@*�LF849��FL�!ݦF�gQ���[�@{W��i,��������{����:��Y�F3dd���(Q�F�����iMU|E22+
��&c��r�e"6���L�w=1ыw�hE���^N�lpX	�M@�h�6+P� ����$�ҹe8���Ȩ��r���_�X�xg���~����$�V*$&���{��	��B�ĕ��"�պ�/�zI]��F���dc7�B���D�6�U�~*��aJ\ᅳ6"U�W?z�>G��]���+�� 4a$�^`�f��!��
D�	(��%C�F��-K}�a��8�c�Z*�
�F6)����v ����ڪ�$�̵Ea{(>�[
I��{f�D҂jV� g˯*�C'	J@2{����j�'�{V勗�8���{�@���{�PI{�_kڈ�g$�\Cq"!�Y�+Q'�����^E+�0mO8g�����`ք~�Be�of��Pίs3,R�FB��w+�?~�GW�uYņ����_�<g�d�ڢW������!��� s���E���FRB�}O�#�t7��T_�/���u�O�(/0����0֞�m���I���On�uF�C|��-�63��O �]G��J眭��%���S�B�`[);OA�[��Gr���	���4�~�fcҪ�z�@�����ð�N��1\�pS���)g�(l�w�'��@Ҫ�|6�@o��T���ޣF<`f�*>�v+!����-�}]�X&�6�.����>��Ss�b0Z(�s�C�<�A�\2�xt(�?���3��/�������[�u\"�����>�v�x*i��9DS�}�2��5�Z�l���eˋ��	H�Rݛ������T1ч���ޡn��='�
Vjii�_w��sf�]�9�4��$Y��I�P��E�*�����L�ǘm|�D#��O=�|��ƊŒ�p�ʎ̔o<��a���/wg��
�Vv<4��ҦU M~a�HQ ����-#��k�H�c���O_%xS_L^��<��(� �2j�'���Wh���+Cj��RwVE���UF�����$ĺ��e�^H�χG��]�}X�ٺ�B����$ũ�D/$�w����kr�K(� 6:6k a:7V��w�Ǚ�/Bb!���o�U@	O�ih~l�L�P�,�������U����+��8 e�nV��KTe��Ş@>��׫W�q���u���^�?:q��6����E(�U�zV�7��?iɑ�z��S>�b�lP B9���v���.�
�M�i��ga^W�_�EE}�Ϥ;2F�npI*h��#� b?�Z��\�I�,�Ȑ27)��.�� ��OMMU	�|�T߽g̊U�����>$."M0��1�HBO��tw��h2h)���'}�cU�]�D��( &����xP���(�9a���[�^�}k��G�)�f�e�y��@@���������"����>��p��n��c�ފ��Q6n�
���@4�I#W���M�'z��4at#�M�e�-�]c��f�)�]�>�F�'�U��2���ߞxzcq�:��&F��zM�%�Q�,>L>���t�=Ú�h� /���A�n�kQ���%��������яf�K�spp[k T� �J�����߼��m=���R R��T�����b�R�9�[��9��!�Zʜ�L̊5��b�'�"O�,Yڥ�*w>9/�F.��%�;��bײ��+ew6K����h�h {A
�H�P�.̧��ɞ����L�)���b�%�d&��!&�E�{�\�c ���Bģ/�� �{�wD��=�_��g~*�-�1h����x9t~��VJ�we���e�������χ����N�����I��b��ч��
��?�����H��n�6'�4����M�1�r���C��z�l�1���P�a�@��v�و\�,�-�gƸ��̩,=(+P��"����]+$P̓��5���5)�}�G��1;�Y��8�e֤s@@@9��$Y�,:��C-�KlOg=g��������5㚼'�+����vχ����p��¬�<���1ǖp#���^��U6%6b��I��K��-m���HHX{���u�a��s����T��́J��_)S��d�H���',����H��{���a��= >0l)���36������1`L`��zff�rOZM���H[K�� �[_0�%�6m� `r��G��w�6�Y�5�y�(�@�~�+�hU�ْ2+s$*���a�~�ϑ�g�P5����������9��f>����Pס
T�n
X�Wc���:Óݑ]9�M����4h���E�U���c`* ��Lor��L��P8��v��׺��1(�A��(Q}OL8JN
@�6/�AjO:{�$Bٌ>|�� �w�G�5+ٺK�b��,u?���,<�Mc�&/��H���XxT�{/\\�=��^=�iB��D� o�]��Ν����)-���C(�Mv�?�-�����o������$�L~�|��_���	�yֱm=V !\?w��q�Uk|��g�@�_�;�F{v �Ü��������&v�o�$VC�a�c�
6���e)'+���{	C9{�D��/�#_n'v�Q��9@I�~��O<�^4*n������3���ZF�>����8���vA�tg�K��7̕��>'��Q��m`"B,U4�L"6���߭�t���b7GE��u?�fŗ��#跴gtT
��G�Lf�|$�f��=�v��f`���H�{�n�ݿ# �ڼ=���l�`^L�
c�p�y*?�0A$���	N%|4X4��@�TR7(w,�W�ZS�SG�boq�&��������Z��3Տ	AK�MeR�{��l��@��	*)oWT@kN�f�A���s����;/�nOz�,�T�Ϣ�����R7�i/�5�8W�T{�.2��f��Z5$h�T糮q��|2Zt��Fk`��31�� ��!�S+���
��92��X��f�.{Z/":������k�J�m:E����T)��$�,~I ��aL�S�,��H��q���"$�c`*���q*?:5���lj��n�~
6�˺�]�J�鳌�HSF
Y??ti4�cR�L�&�;�N���L`�sy��fzo��i�]{^�߾�R�ō s��O��:�[@e�=һ�%�@'���1���-jmH�z�O�� �f��ӫ+�ޝmII%6�9a��b�O`+��|}��g��k�;8	s�>����|��@��q�10r��	�PW�n�x?�#�*I���uT�kdk3-��5I߉d	��NʆpI��]+&P��\�_�k���w�Sݾqَ�MBH�#��J�����c�coB�>Q�doeٛ��y?=��}�ϧ��T��w���^�}]����JaA�K
��7���8��R��3Lo�GX,��*�4�V1h���>��⚣�D*&r�]��1A�&�i$2c�y��Cw��ܡ{n�7h����=���b���O� ����tʩv��/��G6SD�Џ��4��:���\'m������fI�:���+��q%��1ד�6V})D=�v��g.�.[�L�r:S ^���`_)����+���v�g�f�F�ZE�OJ�x5�Ġ3O���pxE3�G�=�<&q���f�2l��6���k�PYjX�`���{vv6�L����΂�6JB���[���m|Z=��^��g�ba՝v��)o��s��h���Dy���@R�d\c���3����CH���]�Pw�Ӯ3��ո�1e8�2ep|4sJ�ܙ��g�_�gV��-Y�ް��>�b���rtk51����wc�>U ����@������E
���R1�A�U(���
S�Q;]&�>(s��P���^���_�G4��Q�޲��+�
t��k9�ѹ��3�@M t������B��zABI�i����؎�gE��}�^GҦ�<�$��6��L|�?D�C��������e�M�-�4<��س�l�P��Mdz�$�"�>m��ZM{�ҿ���գ��ZB����MݥV�t��c����# AdeV�/��>'GgV�!9U�Џ���_b���O�I�����,�-ש��<���9�S�zҝ+��31�.cK�)�Lѣ��ؓ���r�`7)@q�Aó�X �M	����m��5� �P�(AX@�]�.s���<n�0m���i�'��;�K����%&<t4b��&C���9��b3�=���
�@M�4���,io�"�I����&I�{�Yb7��z�����LDE�{�X�V( :�lw�_����p�n���8"+x7�9�l�O�_��G�$�]�e|O�+��ѱ���Z��~Vϓ��K�~9ܰW��sy޿���Wi�n��뺍�VF<�BAfQ�I�`� P���_��G� � ���'��:�~�w`�[��j ���o�<w�?��|p��]�g	)��a\���;�\�̬Fz2)��J�X�W=F.[����GC�p~��V7�M�UqN���:��~iL��1qQ�b~�da�d�f.��U_�N
�Jլ �D���܄Q�,��i}��v:؂LX	�SE��c�v���Z���E$Cj~禜E:5��?7[��D
f��[\4�m���ggd�{B ��.�.5�.!6`�x�B)��
lK.'���Ӷe�&�.ҋ<Ծ�Y�W����`)�nӈu�Ӡ*nfэ�J������G<F%j({Df�?}@�����A����H)_-���0G��B�C�j���2��}>�,1\�3�\�neW�SG[L�d����(�aÜ��<��r�'k����Z:���2)W�_�ɏ�U��uj��/���ͼvva<2x�8�b�/�`M3��[⧲���V�.7�W��[�	F�Cc�SfiqV�7�/��0{v���OPg��[��<��eَ7%8��9��s�}>5�5ꚁ� �-��o�ޖ�D�d��b���X��,��ky��.��Ƀ;傂K��8H2�����C��	���G P�p0�
�T��N�:���+q�gyGiz�oFI 1.԰�õΏn���o�
nΉ�2GU�[pR��)���/�WQ ��	Q��jk4T[����t�a�����0�p�E����{���)��E�f4r`] ���A�	��+��]�Z�EDlO؂��?/~�b�yw�7��e�g�qg'!�O ���f:��Ny�7�+���Y���l5L��wB���,�,i>^<"'�����p߱�R�i��T�D���X	�.����Z ��􌐹�¿%a��ߥc <;,�o{� Xͼ��bN��
�Ut��.�nh�@�Z����'�)�9���am�� �H��ERap-DP�����"�q�c����;Z��[���q��d�5{
R�pa��V�I�`I5eY=U}���1��O-A�cz�`潄��)�[=^��c},�	�1ؖ��,�,^��}����r`���U�E|o1#~6ر!�Ez|(I�kMqp�T�����Ĭ�� "
{�o�_`��Q�S�_w/���f�'���PhjMSK���[�U�+G#�i��iTx^>}�i"(!�+ǃ%�	B��|[q��::����y,�b�cyO<�?�G`K��ٹ�o�{N�Z��F�����T ƻ�NJ"�wz�bc!�Jp�����=�s[���:i{��@!�_)�9�t�
�y
�=��gX�n�_���5?�Cb>����`��� 2}���Iu�Ռe�Ͳ��+�&�8 ��ɼ.�Υl	���C�I&G��p�vi�8-X]��S�x\�l�?�M�sP(d�d� �� G7����b� ?>�_�v��{G���I'��
�5�7 A��µ��yr�(�ɸ�����{}��?Yl���zm�!	�%�Z6Y<FZ��{+B�+���� �<g��*�\��* o�?ۃ�A �Q�� q��`����o�k4���%�-� _ w��r/A�����/4�C�����Qv��<��g?��Xr�·l@.ʀO?x��V7p�V�m��gnzr`ii1Wh��83ή��F܀��J����{������`7�s
A�-���2�`����LM˃u嘋��&�2�Y�;����$1�Բr��ce����f���1�x�:����X����u�U"Y�H����=�G����gI3\*X�1�8ԏ�F͹or���Z~� 9�Ē��7}=	�w��ܳ��q���e�[�{[�^\��w���̤����uP7I�!|YCxr�}�ed�����N����f�K��VG��*�ׄ�U�ܒ��'�Es{Y������Z���O�u�HS��G��DЃ��D��~�)}h��o�ǏM˚%�p'�̥oz�yo����P1CB���6�F1�����Β�a@|D|`��N�u<; {��6?Izp�Y��������ɯ�:�m�H�
��:�M@�>5�|��1saܥ>�u�CW�������!��Qҿ;[=��#���������r�O����d�҄��eὺ��%?!��z��=��_��v9�r�n�?���9�稫4��"	00�TC�D��~���xw�O/��n�I���$
���-IR�G�����'uvR�[B����e���J��w�Q������$�c�q����1N�y3J�CX��(vō�p%ː�P3��;�7����1H�͠��h�������)~�/ڡNimIK��Wؚ���ś���׿?p7�Ϙ�٭`0�)�nA�C�q���2m�wڹ�x`�]Cg^����R5)���K�F׷��Wb��`G_��&���Ȕ��6d��}��\x�	�>c1������$���	�VPLʁ�O��;E� �떛����q���4ݞe��WN��]��"<�@�M[*:�Z�U*ܳ(��h.�����>�m�(ś��p�DI�
iw_���/��ݪ�4�)d-]�0t��k�{���J���T�.�+�$���o�_,����\{�\,󽥖�o� �hs bhUh}������U����E��h�ػg�{1�@�{��A��!rvO��f;�����L�o���.8[�����#x��D:a���i�bmo�"�{|B�IWw�Z��ߪK���\��M/���~}`GJ8,峺���Nɯ2d5h���7���U��M��M,5ׄ
W|��=#��z�^grl!��Ppɳ��NJ��U��r�I˧�[.��4�Jb-��0rcr��E�h�zVd�ԁ������B�g���.8j�If4D��O�*Y;�45�G�1N��r������:��6����08Ŋ��\�C'}�E Ywt7���x���3H��>������ ���X�?M7�J�"�(��M|������}T��ߣ���P�ߺ��[f#��H�^
٫c���� 홮�rR���v\�;t�N�Tf$�w�Rx97�~��/-���"�1��g�]�AfUPEEP(cAD�uw�
�5�>�嶡C"$�ǰgd?�:�>�1�RXe��"����ht���,��:�sP��V������{����?��R�V �}�h���q�/!��UQ66+6��)v�FT>2��a!�!�eFz;0��}.x� n�Ƶ���-��H9v�цu�Q�?a��0J�)����iu!�+#(L����чv����F��kE��B7~�C�M�/)D��
J%f�����$����Z�E�0'�0DТ�T�<�Q���I�����,d�ѯN}W�E�gƙt?R8�ȇvN��N���o�F�C	�4��VGaAu�w�}Y��M/WL�_?Dl�-��n�↸7"��I�,@�e���
�@G �[�G�V1N]������ֶט�c��}j~o�G�>�R���=��'��\�=�z�Y�ݢ"P��9�_��}}��\t��FgҿC*��CD�"�w(� $��,r �\wTn����A$�߻4%&|�h����.��������H����1��ꜟW&�)�l��F"1�?ͨ^�hr\��o�O�ɱ���� W���G���I�-�$+�#��4=�;3wVz��rl��Ԭ%��6�$d�la%-�ճ�x�,q�sgZHN�'QU�4�O��d��@�C���':��X�8����d���M�>gd]�v4�r�|�s���V���Z�@e/>X�	hҜ�Y�$�
�e#�>#nx���a���xۏ�<}%W��C�<:�~E��� c� �V�K�u`��V�`����h�N�o���q�Ni/� �Ӈ)�g.�������9�F��M�1���+fOm������z�\}�8&�wV!j��ן�	@��,�to������f�����u243m��9l|�~�|���^����E�
�)�zu1�	˖@vy��׌.?�������{�Dt�~��&��UO< �|�m�D7s���Ͳ�'�[�u��:�6�P*@ֻ��fOA�Gn��h��a+ּn0S��3@wV��@uZ�T~�(�J�UX�vɲEzB�SE�4���;�k6���0������&�r���$��KYNv,㡄���G�%�Zh�Yps������|����D�����_2��+>��W\a�Y�|:�1�>?nR����J�%1t2�Y6T��*���ϑ�Y�'�$���W�h��"�n����D���WUg����X��<�p���>�q<7�I��Va�����g<?���+��\���'��h�q��n{��`�Z���v�de�� ��w?�B�J�&Qe���؛��V�#(�3���.���(W�Ќ վ$��5\g(�X���^�wCz���`���TxR�A.^� ���o�-Б+��1�%6?Fܪq,C;��q#��i6�:�I�8r�c0PMf9��7�q^���%���Q1T�>�I!���A���� �E�A�O^��!�i�pP�ww�۷�N�`"��ƪ�u$1��`ɂ�� ���<��	�<��9�wQ��H)�<m�0�uZY��~_������8�p�m�)*ä́y��	�r:	�F/"�lT$�5N���U��ͦm�m��d�ю˟������6���x�kb�X��1��{���"��
�o�:	�S�W��8�[9��̅���{�x�A(5fh�%W�$9��>Z��b`}AÇe�d�f������4�Z*��y���_)`�8�=�{$��&ҷ�Ry���y���
y"�z,9�KSS 9(gUμJo�֡bHhE[!���ۿ1T�Q�;
��(�A5wŬǟ���8Su�EO��k�a<��My�_C����d�qz����n�q0`M(�#�a[�3*Id��V�;��������TUY�fR=���e��-�o���[��tE�g����[2��za�ߝ��oUƳ�S�I��<_%�Ɇxn����MHQ�yϔ�U���B٣R�<^�aIg�^^�����)!&��	�����[-yQ���}kC���H��?2P��ц��4;���<���a7 �ϡb�S�Q�f�t��^�+����������m�eW�+�slث�f"m�9QҦ�%}/�s����!]h �p��+_a�M����^��nȣ��1KF�(<�?�^Ƈkm�����_ȴ�S��OB�>���x��W�(ru��:�����6�Gtv�@��Y&�8��gxC��Eo�Qp�		=��+������-�J��Ԗ�
<��6��u�V?mߴh5��𖂤�u�ߵA?{�g��g�R��F�P�Ӻ�u$#�ʋ�Q��|x鯮Y#v+|�J��W���"� ��k����9M����$��M��z��)�'y�P� �D�WF]$1�R�u�~*o�5E�7�9�������16M����ݡdN�%�0��'f�e�MKew�c��h��3��� z���2�f ҧ��e�%[N����`�k��b�З��D�(�Py�2E��	=Nng"�Qh		��N?'%�y]��_XXն��Q��z��VfH�{�$����#�ɋ��8e��\���^d ���u�s\.�����D��>�]�`5�MJ�
�i�~��&NT+Jpn� ��H$`�r,��ȏ��B���j�����t�Wqt㥐�:O��M�J�� �_�n2��ɷ�E��P�;�~�B8�ه���ܩ��o��;x�7=r�8��s��2��� �&��ǰN�N[`����k�=�Z��T@����ӁJ*��o�z�m�U-(��ǵ���Y�Ť;�c�Onnb��G�K��5E��<�p���Q��s}ʔ�
>��E���`�d��Ҕ������R)e4F���V$F�S̞(�'%�c�^p�Q��ˆ+���il��ǧz�ȼ�2������d"b���Z�;���X�T6BA����!
 �<譂�'Q�ؐ"�	���'��!O����ށ!�	�ח���o���"�PT� ls�57��&�Mbo�����_<��Ws�Jb�e�)�jK2S��n��o�Y��M�_����2m`�C��}��'��Ұ}�*�İ�p��z �d��@m�\�,N�*笮�F��P�,N����4�c������ĶVY���_���c�ŶJ���_緦�T�e�U@�t.�����e�������${ћ�d�����+�ѯ3/�b�#0\���6��e,[#.�#�ǩ`��-lĞe�fc��M���8�z�'�l����4�-��$�ಜW�KTO��b�G\<`�R�G`�BO�K��+��0�ǌ����o	eKs0�Е��SΟ,���K笎�<�J�)��� �8t$b��~�Tܿ����]���]�\�=����Y��n|j����]��A�$hn��􎚉2myl�2Z�qk����Im��K���l��g)e�Y��.��u�f��o�����s-�XC����[B��a��ʒ�Ǟ���3V9@V^��.R�e0*���T�W�w��d���۫������?�$l��VZN> �S�y�߿��ޏtj�n�b�'m���=�4�﬛p�����N�'�tK��/ȝ��!u׫T�否�N� ������Go��2V3[?�K+j���;����sj6Spl��G���ł(���)˃r���Z�&S�P\Oq��]h" �*�L��~D�j��1�}
+���@d�g��8�
A}�~֖FWnyM��@��_8�9��
3�ɘ�� B3�Xm�Q�w�y>�Hܒc�jp.M�wx�_�-2(mx�5X���1@�
�s�3&�?��nVc���u8�T�"�Ս��Mߚ��@R�1�Q�hW��N� W�)��"��V|K�����&���׫XZd.���U�~���r�ܲ�md`w�|�_�Q\s2ݨg���2�]}�eCM�m���ץ�5��,�KA5�o������iA�RL5�H�>I�'i��1 b�_b������Ბ�Y0�����Z��O�Ȁ�_������@rF0?P�9���}gC9'7@�'}�4`��Z�
��� �迎2��l�8��F:����"Q5{۝YR�c�))/.K��i�4i4��*�^�lx��-=M|ձGi1k1�:sD�zi 뙅��_6.+�eI�J�H@ch��s�.=�h���U��.�#@�1�ϲ/�d�
d�vFͮ�M�7���IN�����g�'>v���
P�ķ|EG�:`��+�C�1����I���|mE�p�W��h�/����eߴ{��������'��4�wX*��
�+g�N��S%vž�]�wWM9�\ ����`�A@����_����* �����,��~I]x�}��e`��)�qdf"6F�ғ�����M���"N�]�j����h'����O&�g��������ƫ~�٢�Q��HN�c+OJ�PT�p~�c��i�
�v<X?����<`��;e��Q�P���A��ѩ��G����)ix�p�sؠdi��VYc  y%������!�����Œ�/nEBMr�yQ ),��9�Ĝ�MҪ�<`��mB��Y�!x*�֓�U]�Rܟ��.8>�&G]�Dڎ�E7�#=�/O�<�]9ɽ^�`��� p�տA庿��S�#�����Fz�S�[RG��0Ee�A���ɷq��9���д�/��� ��3���΁
�|+�ǩm��J�0Q�V�����&��|<A����.�E��T��N#J�0�����Uazw�%贓�$5��Q��l�Ck��*���,!V㭴�ٖ�ד:1v$+�C�Q�g��Ѐ �_���N��ٴ���m�_�X����Z�  %��<��P�� �,����!�Bp�?�8)]�CC\s�ނ)�ߴ�BlT��M'�0���� ;Ў"'����o�A\c��u֨��^�u*sW��0�ߐ�ʨ�G|E����X<WQ���?��rԥ�F&5ԆG{�>=�Ꝫ9���z��h�<ZM���hC?M����R_��(3+c�����5iJdZ \K66鬊�@��yT
-��wԍ�e w�F{��G;$\x�ĳ��0_����!�͵����&�_Ur?IP8�N4tn��eV,�y<>X���Z�a~����c��"��d�H$w��~��YQ���}@�6Wˢ}:.�?�1�YH�;�fA��oö�pf�|��*�5b�#�C[k�(�:Vx���)�$֝������É9���Ç��M.��ڠ���3�\�k�,���416��͖�N|B}`j��x����%��Y����p��W��������˺d��G���p�Ez��f#���Zt�����Z�7|�o�C\ 7�,Ǐ�	��x'}&D�Zs~�#y�%B��f-+�;N�e���3�^=񹉿U��ۃ���U&��LƋ���ӫ��{�����W����8�*@��B?��w}����%�`~z�K��t/Pua�O��j�q�����bk^AJ�J��R���_���hfw���D�F"Ӄ@�JRU.J���=z=���f�Ƹ��(�eO�i��Ǖ�߳�S�?�6c?wÏ���v��]�<P��곉y�QM��O$���? ;��5'l�����(�|Et�ǝ��l�n�o	#�hT�:�(�1��܍g���]ou�|��Q9br�Z0�~����N�瞔��eۯE<r��%y �;2%��`Ū��G;��Ә�Ĳ(���\���h;�_���.th$~�f`Z��8�u$�#����7��>ɑDs�U�u��>�1i`�<����N\e��1LpE{.(U�n�0��5o^��]�AW1)�vz�CEW��`�ٿ��:}q ]��kR~��T���͈���H�� ]۫R[e����d�+Jf_���8@�1��5$g��
��PW�L~8���/�w���XsP�"D��~�~L��I���ԫg�ILI�J߱7=vJLl]�lG�׶v���)|#[�NJR6g��F���ύV��1`;V�l� �9k�ۤ�y5��=�����i|���mrUb��cT�I�,o�D����ޔ��%b �^�b�뜑���>N���v� �7>�:�ש� �*�rD�(�Q��/%v�XI\g��X��e�Ը̵�>>��Bh��L�~�pX���%�9�9���U���Fy �8?��-OH�W.���g����+2��F��%��<��,���%�LI�r�qz!<(�Ҩ"�숮��s�@d'�p$�j﮼˔��<���5����w�Hֳu��p�fb��^��>��i����z��p+��ᇑ^�?�|�V2�a9)"�و����ܳEtucb�:ŝz2�Z�4loH��f�av׌��M��QޟB��^m�U��1o��h]LʄY���r�K��³l���H�����v��Xz/�p>+��Y����O�<�8�yQ��ւ�H��G�P�M�ռiUn/M�2�h�em�¸�Gv�J:~�7�p�8��!���ug;���q0mW��V��ik��_[;bv6��\�Q���٭��/�I>Q�(��(B�ܪ�l`�����Ժ�$x�%�����-��^aiҰb�������U�6�dG�bκ���fg)q>��%Xԯ���}�Sa�-�J�Q	��X�Rk���<+�i�6�,��ܥ���@�fq3u��F:�֠�m�t�DЊ ����>f�V����ߊ�:�+M�q�g-�.:=�h�)����u-�r��\��=��=iܙ��f��\�{r"��/i̶�B\ɹ�CD�Tf��,�v�����B�� �g����Z�?��u`q+{�<�je��U
��a�H�3,aU�s*�
�䔂�[�#S�Y�˭����E�QVI��]ِ9+�4���@���N�>��yqP�))�>��A�<�8.9���X���[��:�~t�j߳d���)���ʜ!z�C/P�e�[+?��̬�������6��%w/J�xw��-�ƪ5�������`�L~)���)ީ'����F�Ӂg�)/�,n�h��O�O]�fW1���k�8�-�|��H��3a�uއ,k]a����*V����{�|C�7^.�����w%?�I�I�5�(�JM��8d�>��l�?���(�٭�3�r��T�uşŌ�޸O�V���<����]vYԮ�L�\��)u9!k���|�ʩ�|x�t@�)���6/�>-%���#��5f0���=4$g6�|��+j��zkY�"���l�Ft�(�ڢ��d���O�R�*���Fr���kqi�F1��%[�Y���'l�zd���S]�o�#��}��yp���s�g�_�o[~���F���K��'��V*�%\�� ��˩6g�((��3�(�����m���n�'JIܾ}3��#��y�V�Ǘ����f	W'+˘�muU��ӑ7�����`iJC���\[��X�u?F2|m�2`�@x�p&���F��B���8 ��C$_΢Y�l�������l����M��&>�|靴z��Rgi�ɯ�_ �H�Bn�s�l��7]п1*���>b=����a�y��NE������2�'�p]W�����3�5�7���Әá��{h=�_H�6c�Vç�7�&�E7����
��α3��i��R�Z����`;6	-�̹�B1W����a����%��ϑ����s�0�_�k��m��a�����e�8�R�2���D�|��`�OWl�÷W�4��Q.dYL��_��y�_��p�z�-�^ִ)��銹n-a���&�͆��}�y�B��=��cڄϰT��N��Zݗ?��s%����3�h �P��'�X�ٜYvO)v�f뛹�Op;sb���&v�����X�Мd"�Zo���~��mo���V�G;֤;�Ȧ-�󽷰f���()�^�����lX$J%Ir*ۆ�oWOm	@��&�+UAf�̤K��}c�;5�y�v_�9�y��g�ˋCl�+�_��q��- =��>�˨�<O�d|gk3Z����^�/G�b�a�eϒ�f�i;�v���c�o`�蔍1��^?,��|��O8�d��ſ�E����a��m������� �Q��ˬ%�nQ����nM�T_)��`Y�h�E�ꛧH���	Ꝺ�-�N� �!��O3��l�GF[�{d���\ξ�;ԟ��3�3hϕ �
�i�����X�5�{�e9��l�(�b6���Ǹ��f9-W���KdH}�Y�R���Tx�L!�X��gJ��,��0h���ز	��Y��"��,�箱�M����X��i�t�?�����_&\G�����V�������x�;��iU���PK��oVH8;�3r.ȝN8=g-���=�h;���bA�}����4?��{����n��E*��C�"ނ��'��q��6)wR�(/H��r��h�f5v���- o�Ua�4�D Z|�"��_*+�6v��2Z2�H��"���n�u�}�/=d-n�����7��A�� �&S��]eS��}fW:�$�?B���~p�f��%%�~YBM����x{�zp-Z����3�Q�"�j���}��;#6�pSO.s�f�%T�G���	�(�b�HjoP����G&_^Y�!�î�ehct-���U�����w���r$�����<@��l��d��Ҝߣ��gp(��&+0.�����}���3p-d�Қ(��ش'�]����wW�vaPwV.JDO<���$��D��n0Y���0K������fEgZ���5�z���������h�B�l������`[uid`Z�+�̖)R����0��/���6�L7��g�ɡ����u�>yh{��D
�O�Άb���ʆu�^j�����P�ƕ5��X6��ٽl�#a��ߐ��(+(]����V]m8��g���Jb�֕����&T���JZ�Q��Hk���0q]���b�Woʿ�6��ach�2�4�n���ɵ-�zW��+�b������ңg/M��gn3C>����ػ�KB�\�4�K�ZSI�Ӵ����W q%-�U_��|���V��w�0�"�>��.YSw�[�����Y`ףF-4 �X�rx�5�_��OV��4��<��	�2V���+�!�2��VC�C�0�x�OKk�8H0���
&T�+F�HP���J0�R��2>�{B8�G�g�.���ih���w% 0�㉽b8U=�y7�R�/��c��,G¢v��� ��*.9�:�$Ė^�����JO���Փ	�嬋����������cG�31x_�""�
�V���{p����J"}��y���#�J��|f�%�͵���qIɨs*Վ�'��1\���!�_`��~5�aܷ���l.�?s/bq�]�l�S[l�B��2hz��j"5���@�Ȧ!\<O�/eWy�L�y
���S^�h-�2C�(u:~<49Ho����������MƊ\�*��∽��ɚ\n�E����a*.����s����jT}�n����I�H����/B� ��Eb�<Xpʲۻf!^s�6��Xa�.�5i�m}�=�#��7�G0s�G�۝,�o���	��~O���d(��9Gzsd]���,|������A� �&T�`=ŉq|F��0����^��s��8�L���Z��jx|�ջ��^W-ah��3F�����]{�@7��DS+Z}d�����\�A���)l&���\Pm3WaC���y�]n��ô0��k=E��t�*Z"��
��_�/�߯/�6p�
�?�q�����VZ�����;�����<�Z��{] �����Q@�L�G�(�~z���'�\d�B��7���~(�B/�r��S�_F���t�m�^5�N�qG}�l �~����OD�c������KϬ6_��YO��j� ���]��P
�(���8&���5u������r(������J�[�U2X�����(��$�Kk^�W:`������Ko~�����T��X ��3��;G"�%�B��3����]��m���Ŕ3;�-GVN���=2m��V�;�y7H��Z�Yf�:c!~���Dl��a���(��#κz��X�����*�_����K�j��1q��h��&�`t�̛s6}a�g6�>�|ƿ1$,��ﲒU^R��@De���|f���<t3�@Q(z<t7c"ߥU�P�,C�[D��wDE�-�f���#j��?=��c~�*>��'H��մ��������-d=�Kh!ns��#�C<�Aͯ��*�S=�����J�AO7�틟��S1�ߺE��o��{ݬء�ĥ4�� ���|�1��߷Vf��c� �#���D$���g��/�֦@�=�k��ս���i��#4�\w7��O�(���q����9Y��#�w�z�
��NS?���6��kY9�:�u%���]�ͬđ�a��֥�ͽ��$c��������;E:J�gM�ֵ:K8�����c�smD]��^��x�w�?�$����j���[�N�׀�H�v�e��E?GT��F��2�����������@���b�s*��\>����������wg(��=�&	��j�v�a"8�C��7�M���`@�Z�b�)�)�����ޒ� p#��(�������ebګ�}��w4�C�CT$�u��w�{��&��Ubr�8Ϋ�����g��6���>���A 8�̅D��<��������ǆ����)��¦a����3*.W����?��u�3����m	������-�d`_��%����/��������I��O�.�%-�h�Q�kE`1�"N�R.q^�R�3XQ�F؎zA�2��WUb'06_��i���8���C�5���8���
����RX��p���L�D�y�Qx��
�����.�h!9%W
z�jN L߀��w�~M������9	��a���8�?g�>Bq<C���	�]ɅM����Z1 �N�g]���3��s�:��#�?�l,u����lc����H�	��!��U5�hy�E�ޘ�wĺ?�H�c��
�j.�2H0E,T^IyR
&�����+s�E�f�V֮��(Gv#TG���>q����6
V8pZί��4�� "�ai�:��*�@��˔�WK���d�����ɳa�Y8!�nApx�t�t��ǿ '���8I�I���Ν�9_^	<;�3�'���Ւ����b������̾?�Zb�>:Ϟ��1���J��j8tOx^Q����,]b��������B���������ah/���nk���W9���=W��B�@u[�~	�bF=!q`X)'Z��$���,��.,b�j�?��_�v*2s��Q�pp�i\��{5��ef�V�'n�oχ�����zq��Iy8ĸi>�`�bׄ���茱��qȐq�d�S�xBh́������w�xYÒ~�r=+�nC/�QϮY�ewϮ<�p$_/`���ݑx��n�{X�1�:"/�!��|@��p[��@��g���P�T��S <��b��(���h�	�0|�,����� ����:��E�����lM�5�"��뱢[Eˡ�	�R8��?���X�Ã���Y�|�p���~&�f��2��;����]��otv��'Ѭ	�Fa�������%#b��pW�Q��S�WP���k}������?��9�i�hk���G8��I���z�z (�0\�˃@nJ�h���v����ME'�;�N�L����eo�n ���E��*?D�~� !A�G�q<Bi�2YY0H"fb�u>Ѯ���s=��j�>�"�,| �A���t�x�ڈ��W�J̎��a�,{�5?(���c��m���?��(
(�)A�>���3�ޡo�}f=�E��*$�7+7�4CINZ�+���$KkXt��F����F"�rV�ߣ|�=�� �yŁz�B�Y�z���y���J�xD�����y�16�[)�r��m�D��I.��o���M�s@C�P��[�M�
�:%h*�!�����iv��FG738r��n=��O��Gq�TNG R�!��ns�7���S�?Z�}k_�żXRl|s���p��J/�Ϟ����N�uq?zۊM��[��+
�\.ڽx�s&�U�����5�_��d,�
��yEy����#Z�b�=gd�Z��9%�%��8��Q��ۏQ'�����9���5�H og.��;�������+ԣ�X�~�I8�Hhh����s ��n���d<b��xܺԓЫ�Rc����_��ڍe�3����YaZ�2��$i�y�O���*�ܴ/Os��%�M�1
�?�gU�S���h�h�:���(�x��MA(�7�W�ݻW����x!'p�� �f{��ֺt�N�ްQ�T΍�װ�ڜH0���d�9��-kX+kv�͸�S�a�q4�0����?X�D�d�>*{9$�� 8���k�0"N��|�Rj�oC���F㢊��`�B�Bc�"n�����Ew���F�d�.�Vn���3��O)A�>D:=�}�7Vn�RC�k"���M�t����>~H�&:R�\O&Im�ˤ��zN9����o�>BBj�4�q�wL���
RTϨ�ylv�t�Y
�ҽ�I7����#~%j�s�1�|S�\��T@p"�7k7^�NP�AC5��3	=�,�k���� ��>���5*������x�ɜWT�T�LM{i����M����*�ݴ�f�#��~  U��V��+�|��h㛟vշ{Pt�w`]e�B:'�RJ�� ˠ���0Ŀ�<q6������_��vޣ�崢r>�P��"ɹ6�2�+�4�~��Ɂ�V6O�|��?�}��YHz��	~Y��
�VY7�L�C������J�$le~^5q�1A��|ʸz�sv��Z��R�Ą��"YA�6.��J���C�PF|=�w�
��|8ݙп9�1T����	��vz@ø"xz/�<B.	[T�&�I*� ;q��:��$ҋ����4������tx=Z�>��������nM��܁t��m���He�#���l<��X�H$�I�L��b���+�S/`��I��)CE��F��C�����ʑ3���IAP
Aפ����˯�	~j3oT[ �;aH$�hZ��C[*��eȧ������w?��F���Ї*o�V4hkEkojԪQ+��Z-�I��:x4�V�U{E�Em����V[�=���O���u9׹�����r皞��bfjk�+7a;�R��U����&�Y4{���k�)�x��]Ks��u��]�S�g2 Q�_�}ލ����tu�&+��W3��(R�P0��?7L�\k'N;�ah�%/M{}�m�S����k\w��Sǟ��.�Bh�U�����t��ݣ�������������?�y�/���8i���'+�'zq>+Q�����-L�`�{�I�}S��ۛh�`	�E��٫ܪ2B���Q˺@����%��gj͟�5�K՟��X�R/�`�O!�h6<y��id�|wro_��eX���	{o�!��&��?�B�?��Lo?yT�"WN<��"ކK�&S����'iK�+^���y���I����z.*Z0y���[�Ƙp�Z�~����x�ᏏO^� �h<�o���M����o�r�PA�����}\ �&)H-�K�_f��!4&�ض�Z&�yg�R=}������Cϣ�nƋ���k���T��fmvrc�:���ӗ���/����a/��HH\k��
���%ұ���w��󼪮�%��9Cg,+���هLx�k��_4���M#:�|�.#2Vٖd�9�_��H"n���IFʆ���ы�hp��[�B�Kl�c\�P�<F`x��U�OE�Y� Zh�$iv���d�de��ƃ9�Nż�/ ���1��7����rq�*U�O��w,9l���z�rH���6�ɗY(�O\@'��d��d���e4�v�*8��˄������O�ۣg��U���EC��&��F�fuٮ�m��i<'�#79�y�0PL���O�KB	�%�6��o?<HJ8$��h�_���iF,���s���)���ע_4�k*?c��?���'��K�;�7�kJ[�x
��"4���<�D�z!��^����XC0ݼ!���h�E�sNz�����N���n���!�P��I���a����<�"�2T.�?��kz#3�4�|ۥ{3wvx;��q������nU��B _�,�}:i�z�#��b<�jTQ�Κ5��N��bK��l3bKb������hS�k��W�?��I���C�@ И�XO�}��;���h该�����U�+�q�M�� �z�J�瀩˼=�ܦ�D�>L�v��5�������o��]_ވ&�
��!��`ٝ�We�F���7Iʤ��r/>�&�py��Y��Q� ����}?���j�Q/8����2�
'Oe'��嘵̂&o��=�Sâ:����m�,����P��h�q��g���՗�T����ߔ]�,��\�0]��/Ry�j��ģ������TU���R�`�ǰ���7�j�Ɯ��9\Ƃ���N?x�٧LY5TQ� ��Q�H/�ё~���v�������F|���<�&�+:&�;h� P8��1��i>���������z�dl�|]S^�1vo�����R_JHj:�f��@��4	3m��M���K����\D�¤���Q�}��1������Kʘ�����%蛇��*�l
��U��Ԏ�r9c>����4���ן��.�3�.��&�dVa��r=W��h�+���VX�8���!Ǭ�p���s���-��BƟ��0r'�%�$j��+v����Ji�����:�N��W�kv�Ҥ!U�w��+����k|���~�syk	p��	�+x�(�i��1�&��!��ec���e�[�����$"��h5Cs,9�*(.�6�&��r�vx7���;ڬ�#�`��S�s�����H�ǳPP�W[�6tr��+mt�a�h�� �}Ð�W�+�22i:��u<�\\ҷ&��r�%���gz���}ru�}��ʮp׊�	}��oʉ�|�������|�seI�Mg�{�[g�-����yI@�uO,����w�S���!�
=w��	�Fѭ�+|S�1�7�D�9߃����i܂�T�}��f>���(P7
.������,��U4@.�p�I�`7n���3P�1)�~��9a�%��b�C˴j�FX�叿�1c�/]1	ޱ��4���'%���R�|G(jT��>F�:TQ�4�+p
�a�!O! )ԗHnzF�^�*�ik$�Q["T(���R�b��逽�22]y�{���uE�=|!���ԁ��ϭ$ez�M`t������5M��8?J���O`#C ��q���fޢNqRe��7�Q�6p���R��5�Έ��x�%/��u	
�[k,Ț���x� A���\�y�kG��`�[�P���s�>9u7�ה���j�/�0�\ ,�ny)/J?�dR���£�X��o�H��1�p��<�v��=Z;�m51�� ϖ��[K��|�z��M��pt��Q�U�)����S�(�w^MG��]n���!�3�ΥF	GBC��#��r��Ҽ�f*a�O�;s?]�:=$�o1X�7��6�����CM$�3��]WQ>#`�j�٣~3�= ���ll*�9�?���7<?��쵶X�V�0o�g�Iy~�3]ۃT�� �9h)�N"�F�Qɶ�u�4| ~4��8���;���pDC�t������	�֑u�sY([�ӎ�|�2�����R�*�f�I�qs��fH߾��� %����c����1*�[�`�l����-�(���lKm6���tS5�p
��-����/%̛�z��u���F!��0֙�x����cE>Lb<�A9���HU�e�vIo`W'�v�U���Ti����x�xm�W�"u�?��t�%�KoD��֙���S\�%IoZ��iu�C"�`�����{ǋ�2�ۥ��n����G���v�V��B���eO�S�f�P�,06,
t�_���z'5sAUCzA2'�([�2�D���~�(��e�X��1���M�݅���t��6�z���wX��.�׎��7����X<�~g�T�nѬ_\.~�;��Y�8�ׁ��dكZb9�f���3�1��Ō���F	6��.!�2��A��1j#�>Ok4}LC�~�CX[k�n(���t1�:6�����{�|k�q	��4�b��n��{��/cs��ڻC=�n����VѦ�y������Ȓ�1* �n�W%;T�4>�!�]��2_s�>��ީ�n�pޘ�i�薇s�t�o53�H◆G�F�7C�@��A<1�:Qå��ۅrP�ȩ��8
��Y�'
�����BC��(`e�6�0^�yEx�}#�_�_GE=�6�"A�c�!F=���S�ȜoRsƬJ1j���Q�I@��Ƽ��5��*~�N���G�>Z�۾:V�x���\�N#����}F�)O���0y��k�$�n�L�|��<�}��Z�p���-���2z�����Φ�^!ݦ1�R��0��d� b��ʯ��t�&��Z��Lދ@+k��A����z�]�܈V
���b�꼤��H
�*jMS=:�OG�%,�u7�>�K�'쭖D`��[�5qۋ��n���^�l�0IN��T-��$=���'�[�����x�̷��Ig2�ot,��Il�=�2��m�75�[�j�$}��nx󕘇�Vc\׫gѬT�9Z���:�o	�gY�Vc�x�@�^���?C�����h!�k���T���"�D�O;���@�����{���k�3��ve��h�A���'�� @�IM��~�CƝ.�N�$�>�t��iûY-�w@�Hy�*fn�����n�P�N�;8��s3������5�$-'��hȢ���`�4�gnqt���)7E��R1��k�>=������sy
�X��L1o�4MgO6�;l{�ɍ֩�G4�q�U�'�]�^ɅI��z]�tW��c(q�1*#�-J�&��1��P��[x���ʣ�T�ӵ��[����ͺ���;l:�)�Ʒ�6�8��_GD�<�&�~I�82nk-Jri[��3�D?����ð�&�T?q�zSR��Jܼ�s%�ve����<V�h	�k��ʛ��(&"��OSȅv
{Ü����W���K�!r�~3�.��-ݕ�D[�����XČ�gC����4*<��C�c�xkg�k��N���S��g*�_���eQ�"0]�֖���x)H�HgS�����W�o:���
���%=�Q�s�y�8�����\�K+ᩌ"HB-7��<�I�����kA��$�w�}WפǴ�Y�����Y7_��[�4�a�����`��A���ά\{���m�Q�|ݕ��I�0���폰i���W|��3���F�DݐA�~$~�-��WK`���ֆ��b�'��!8e
i���v[���VZ��>f�'XǙ#�/ᖒ*����Z�o5��8��YK�L�A�гτÈ�uܗ�b;�m"i�΂���;�@m���� m�K���ڳ����K�Ȫ~���T�w�;�S<o1z%�p1.��v��H_dC_�`⥎z�� ��K��U��sF2 �E�`QCն@�H��/��v�	SP�2	�I��S�hM�T[c::�3����D0(�ˍ�W9��Af-�g]�.S6,_�mJ��)�>��-�	��Ujڊ�GM[��.�:l��#�]�!2�k=0�Y�A��c��q�7��{/�&x���|��3���N����©I�ǹ��{¹�-�K�q����}4#25�'-�}�p��׻��ef�CN�T���^΀�����`>w�A3�X�(�� �%n�r�=��صUD��1O�l$��ꊯ��1iަc�?j�8����^X����YUe����Gu*�b������oj7�t��K��ʴ�$s���&������P���ᠥ׭p
�l;�P��������wJ�������G�F�����Um���&�YO�d�2��ۭ0��]@�kS�T0�|���!�ޞ��$�kǍ�B��Qq��&�tE��T0�v^����M�OA|�@�j���ͼ+ySJx�ސt�����>�3>�5�R,�Sn�[:{stH��K�?Z�R�E�h_����X���;��k�u�S�P�����/�f|�,����W�հd˵�1FT������{1ޯ����65�X�G�ps��z�̺����]����q��l�W�3��zL�O�Q@w�7��ɐsC�p���n	�G5�d EG
\=^�`��ƈ��Q��2N��/o��Q��m

�u��3&ű�(%ؒ���s�/ҩ�N/-yVgC�Н������W�wK��FP����Y�Z�,,�2�%����;C�4*ӊ���+2'�G�5�T�� ��W�Դ-�K�,G�ka7h��֌��9fޖ7WߏN �F-g1l�y�{T`�����vٗ%=H?cߏT���� "��\��O�I�+���ݠ�)�f@/�ꁨ@��R+�%q�*ݱ�U�D$�Y���H��L�Y5��W�9f�`]��23D/�ߐ�U�z���=���%����y������b�՛:�M�=�Y)�)�1�%��p�Β���%���{�A��h�����]�����<&��/���d�h�L�zaV+��G/��Q�H����(�3��K��u�A���v�ܕ�9Dڧ�}��_��^�C��<\
���&�HC������I4pX���b�%]H���{^
u�0��g���ԥ9˓��n���X"$�������a(I���8��ţ՗܇�m���[�C��7X�?��A�_��z(��(p@(W�/���`�����L3Ot��I�ŋa~D�1$Ϡ��eS��LꤧKc-u����9<���Y��X	͖�t�[�1wB|��[�bMww�{v��L=I�\������rt���a���J���6�¤�Ul];��ecڣ;�O �F/��ޑ��}��T��ձB�#8�8p���$�!j�-����o�c��.�h�)����У�/J
�>��Am�4�����Y*/$���W����X� ��@x�Yi�߽�b��8e�?�L�!��:��6'��W�Y�~�l����6#^
jfC������R�ͤ^`Y?O���4�������ȑ��*K7��V�h����l���߆ֿX&�rø||h̞:ed�����k���(�ե��Κ��3Q9��[�큍?+_a��0:=d��N�W���#]d�;I���8-9Q�;�I��k�V����_I>��Dڌ��cF���ԳQ��ҟ$kw󺞛�8�:��g��ѵ�6�K$M��V��)+����x��²&�?���7�!��ݥ��Ԣ��$b�$,�Sk��HU`�?����q]�/q�8)|�T@~�P�RU���N�ۍ$�/{�=��`���M��ou�S��i����HZ��rj�j.�={,���� |)�W�򙥶�}M�,���z��Ш�h|;�7	��Zz�ՠ��T<��
U[�N�|�H���~���O�V�a�S&�l�⡬W<#E�!J������s� eb|i�:MF�����8l�q+[k��=G)H9����t{�]pj�~��G�T������ga��j"���ˢƧUO,Nz�2�z-�e�����ħp��煳�1r��_�c��������6	q{	6�s���kMmMrS��	��!=-��PE�w����_C�wܢ2��׮8w�5T�E�gK���z��]�h�¦>����X�W��f`�;���͕}>�Nw[.�	�)���h¯\eIz�{dBۥ��[��O�xE/2;�2Yn}���x�|�x}�I�@��I$;g�7����=����_��J��uW���B����- &^8�	H�ܘw�'����'�,O�HW�9�K��"����|OdM$��Z�EUK��ه��WH%}�������}en_���épW��1]�Cȇ�O��|���P��yB,���q10�&�c}v��9M�UA?����Y�{\���0�N
�d~�|��9�k����p�9�����y��(�s����]Ǵ���E߫�������C醯VL�&��U�����7�,�MHK/�V�/ì�PE�Q��9�X���C����������l�ld��~Uޑ��"䆇���)���	��~�=��Dw%�M�~.0I J=RBH*�GY�o�{��=
��IESu��/���i�&K*JyM���#8&E���[ZPNI{�*m�����@"�4��6�Oi(F����������h�����|_�>�|-Ѱ٨=t��?Y@���@ۣ�
�k\`U�[��?�����_�@�γ ��9�@�������ϗ߰ӹ(t�����2E�|�go�PK   �p1Y�7}b  ]  /   images/cccccfac-78ec-4b9a-a64e-108b6f3d2b7b.png]��PNG

   IHDR   d   3   ai�   	pHYs  N�  N��"��   tEXtSoftware www.inkscape.org��<  �IDATx��\	��Wq����c�{gfgv��5۬/��)F���("�X�+R!"F�����#Aز�m6���]�w�;;;�s��3����w�����O���.�ݖ�7�]��zU��ޫ�^�]���>D��)wb�d�����p8J�M��x�Q��iH�xڇe�3̣��zI��V��ϝX&��\���U�9��:f��h�P���$X�pbf�!oV�+��
h������i&�j�fJ���Q��0��� �97:�bН%)���#F�w����<�%*�V'��z��fs��Qxg:f	��P
5�����i�Iöi���S�o0y�����)�C�����Q��7�{� 3���p��ӄQ�PG�!�U��;�a:�L��	̡�߻�s2�k�2�	�;�����8�eH�<J�Q�"ux�n�`DC&'��`�0\�`�5ޥ@z�, a_V�i�B�=����e����qd|l������E�{:ZW� ��E��{(Ң{��v!f�?Y�������)wsǌ#��q<?�B�%�*����М��B����ᖫV���qz�O�T���L	���&X��^ӖAS��'φ��u5���˵�^�:nqî$��������ݽ	��fI1�M}o��!�v�8�v ����XN�7���1�<�䲻����%0���ଯ���z�486v�3C3��SC!5��jΡ�)�Gτ�1)o���
�}��Q���Od�b�Nʏo`�)�ߦ�eXm�ؘ�.��ߝ$'��F�%�􌏤t=�����6�`��[	�$t"f@��D�If�ҷ���Й��I������^"WXc,!X%�6M#��(��"b�;+�$ac~�c[rK�J���.��?�u�|h38�X��k�R�f���1ˮ�W�c��^Ni&�X.�*نd�K�,AzYU�λK�D�E�
�'=�$uWI/�F�%�ؕ�`)��� ;Bm���:�t������7#}s���D���Ӥ�]�0���ۚ9ƶ��y��ʙbO�g1a��!�b��o�E��I.K+(�ؠ�P�pV"m�M�M�QOjP��2+o��l�4%@ӯ@_�`3�-�dn�k߇���Ͱj���c��H��drVJr4& �t���	�'�u;������Qlܽd���\T�E��P�D#�9�&"��^�	�6U=a��(ڝ��r�Rdx��!���(�</F4j�%�l�g���G��w��[xn��"�V�n�S���,X��1��V�4p���t�&Bv��P�,a��*	n3� �A�4�{�}���y�m�h�#�����(��wt�&Lj,����,����&��6"�/���4�B�p�:[���#3����Cس�C�?ta
��*Zښ���$��S���mGMM~�h`t|K�q�j/�~�&摜]$�;��gjk��,�p��d����#u����1��Z�;��X+}��� �UD��W��u#��`�ܸ_}C#:;��Leqfp��\�����	~�|���R�>�g%���㖲<�2C4|�8�
�Ģ�R%���l��M�%�]�o��d��	��H��Ko�V�5d`]N���ʩ���P���ġ���IֺX,PZ��2Lw�|����@*�&"9*�P���JR����&L����U�A��ԖN�x�j��`�}�v)U��_P�.]G.WRmҏ9T'���ߔ>G��K�_�Z��TFn�p�o�M��ot|Κ� �t*'F������
�h�Q��ф՚��XM��K�Ee�w��9�7=�$�`0�g���<�BmiV��Ό
���C��C�E ��@3��Bx�0>9O�Ε��Y���qJgrg!�2����2S�o�����ĩ��*��R�X���s?���VI�%$��a���vQ�]�Q�l��W~���tn�qc�[����L$�B���-x�bi���� �����N��l ;щELN/m��%1dc*)���'M-��1��b��084����;�N�q��I�����M��>���<�+�&Hsش��%uLل-�V+GL������XZZ�]w���_����'�p:���[m����xu���ɞ�������Z%�����u��O�63���"�m��������ӆ3���'n;�mm�HҶ�c��<r����|5�UV�|m�k�:9!�M/�gf�h�D[��ر��BKf���dd��%���<v6���r��Ѿ��ؠ�B~L�,���w|�3x��1ڳu��u�p���ٶ��,f
;����Rf��[*����,�y��7�=�N݃sS<��������*�F��jIL_�������S�s�\d���=�C��`�LY��>İ�&sCG�_�닸��G������|wC|��{��lY#������S��u̷��3��1C�]�Cf���&Ƹ���?��]�+9��7<C*��$�.�F2M�By��e��/��LF}��9����s�o?�.4ԇ�9��lr�Y?�啛��ێ��%�%Mՙ._U�,�6�ȯg��c�V|ʕSY�T�������(�JkOkR�07V��夻��V�; Q|�t۠�������(��ne�uy�:K~$�����o�:i	g1�⛿�AW�Mi<p��*a��.F�.�ZBg
z��x�/#\X������W/�POL���tgwCڒ���̹_uy�J3�
.�dc����ئU
۔]�)a'.[�����zJ�y��Sg�w�eqxw�4�//���L�d�t�^S�&u���C�꼁w����l�S�P�:����V���|܃唛�*�Huu��S_bWJ�oL��*��ģ���>�V�8�>O�������n��c��ӆ��9!�}��/h��c�rN��li�E׎f?y�޴�ӋXX\�C,���	��I������D"]�������*��thW� a5ľ�;n^�(#��K87�ώ��:� �O3����������o��_�^o�� �M ��������|��9O�L��_�w|���G߇��>bPZ��q�¤����j2#g���`����� O<����0�����<�����u�a2�����MfO�[ɠ��Z���S�g�3r�~����ŗ.���dp䅳��Ղw�z-j�|ph�iF}�� IG{[�̚���i�v2Y�ֆ09� G��\ՅPЏ=�;��{�M7�G��f^A�sYe�g�o�$����h�S7Y����5!>�|�]b+�6̱Cp�������VM��A�0��3���~�� >����} m��8sn���b��S������8���)L.�֫,���R*�Q��b�:1Ad)N�B�ňo؇G�|ѕU\����)Qao��]�z4�u�"���BLȡ���lC1켨���%��.3g��<Bjk�;���݊���T�V]���ZA�/���Gv�3��n��:ë�'|�$:k�djR�=�����f_�x��uV�RM��5�J;l+N�ˌ��3��y�lۈ���Ɍ`f2sy�����I�5��f����u�)�3���o�&vܵw6�=�p�/z�qg��n�^�sn;��XKj���;*�)֗S�e������Z��՗�Nx�{t�5����U�I�����:�d�{�� �E1�LM��e	6_�s_�.���W�L�h���λ������M*]'՜�����ǃ��O�^��
3!�+��<Fj�g�f�`��p�>��>���y��� ���7ϋ�2���5��͠���o	�xjU�d�����u��� �mwh��O�����+���]�;���j�q�����a"�W�Q�R��g���|a�[l�����L}n!Vv�t���k�z$���i�V$2.��mf��VY��Xd�*_T�\m^�jȞ@�&�~&�����m��28;p�--�����S����h)�yѠ���r�U��y+Icf��qo����=Q�U!�Wބ�ZKl�x���ބ��(b�8��owbp` �@ ���Sr�w���jo%��K5��J���ϊ��nI�
�3rE�kz�c]^��$/��Ey/��y11>�CC��|H�i	~��W���Č�]��юK��_cؐwv��ҒB�z%��.�PЇ��y���������;�W�]C����7�n��KM���'�����;W�0艧^Bm����rs��sϡ��7�r���En.^n��b�K�tPn���U�Ea���M��~�-�ު��iټ����M^�b	�������x\�`Ng+��pb�1�NDԫ�-�e<؁�#���'`��m�\N
��3rH�ʤv�k��H����񤱶��v��&5`Xul�z��Y�`��꟫���G�	&/������tխSG�o����m���6e����>�ۉ��4���G�mү�򂊗Y�)�B��+'Fpwo���W�i<w������߅��Z���3Y�85,������\�wp�.q�O�,b|rA}�v�s��%��oO'��=�L���:����?o��}t�h��؜<.�r�!�n/�i��>,���xF^4��r�Į��]��������s�s��ӄ���j���*F��RG��/Z	���=ޗF�u�^d�"��3gǅ��a|��ߧ�[��b�)�Q���(���y���~^eXXYB��Iĭ�|�`���I:�f��+�����D���-={�/,��cZ2�$lq9A,R{%�J*O3o��f��Nb�I��/�^���ȬH3�V�g
>�OpD���.��0F�%-m��T���r<��Ub�z�-�+���g��$p,�[̀{M�E�2�8'��-l3d�	����)�!7R�]�ɁD|	�ļ ����`bb���sI�K�4�#q!�a�h��[o��))ǁ���U���e5妁�H�F(�L@sx�r["6�Ċ������C,�����KF>���*�y���ޟk�o���22Ɉ�a�R��,]�*r!YD<�}����1��>L�1h,��g��D�dB�1ᮤ� �?GDP�+E��H����Vy���R���6n�yЛE{m\�ۨ�.ڿ$J	��9�連)��@$F] %Ag�eeM"�p���`w��8� �)�j���ql���0v�.��l܏�d������.�f��9ڄ��hJ`;ڄو��&8��S4T���`Rpb��,�֗�ߓ�%I``cZ+�E*M�m��J1ֳ�2�8��͕��fH�̢�;�Z�#����q�1b�	qdP�:�!W�Ys�S��80�S6��r�KĔ�Vua.+$�n�@H����J�S�7�'PD�`�DtuH��ƣ>�R�C��� �0��5��T.�х�!�R�M���c1�<u�nn=�Q(2���fB��pq8𘄧AL��Q|�.��7$<��R��M��� a��z�����k�۩�����o�|����l�WgZ�眛�єV����2¤�-�7KOc�.Y�rT9&�N��s�F�2��2��)<p�N��%?�1$��'�T�	�Wc&�N⡗k�-ZoΉ�o#�/�D@�0�����^��-3��p�R�f8�U�9�{_{�F��)���а�9+���p���b`+���ٰ�&�1��ud��S�"�<�0G,�MJt"���@~��^b����jl��J%C>C�����,TȠN�����D��χ�s(��[+�i�d�T���OPqY0V;cKLF��rr�鱁�2�$��	_y���-��,��c*���\PS����G��̡��0�ϯ΅����Ϗ��ݹ�h@چ�G<��S6��YqK@a�5�(1��ӢT��d���OBE`�G���Ǳ!�ɏ,6r���]f��$�ӎ���3D7s�2���G\k%�(G\sav���}������k�f�6����0�;Ov))1�x@���۰:�J���a�r�yC!϶��b�hk �dG���Nd֢ޑ�X*���^�.kE�c��ޱ�d|�g�D�c)ZQ�8��4{,�������L�����a#8�}�t�?��q�d�    IEND�B`�PK   �p1YXs�銙 � /   images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngl�T�m�6<Cw�t�Hݠ�(�(�H�H�HK�tww*#Hw)=4���>�s�k��Z,��c�s���M���2>5  �WUQ� З  �\,�'�~��oh.r�����/�E8�gl' �������.�C*WE}W]GKW����l]>�;}�u�l��� �
��=3�=<���1���/�U�Qq��hZ���DĊ2d��s>�u>EYẼ�SP����L�H:���pt� ;�y�o���P(C ���ȁ��e�$���)Й%vݚ �������f< �٭�=���:*�������0J��	���� Ԙ *@F��u��}$�)IzFf�Y�	��$��;��8d�+9������%F��-լ�u���{إk�o]s���W[�Zx��d�Y�9��$����ʹ��R����a�%燷[�2S������x�9�w;2z6,���2���� H���m�z�#�2"(���	�X�w� �/�q�լi<hk��.��\�X��$O�߉��s�g(�4'eh�j�w����Pښ�ᣔ��'�K�sI�NY7?ι�X^��2����D����/�<2��|�|���F��i�ŅƮ����5�H�Y+u�7	з\��NC�/�����dJ���:�^� z71���'"��gl�n$�n;{��h�t����u��va�"��bEie*�S�c�#m�t${F�滬�k�уQ�9��v��@�MW&~�[��l��Kl7��v�^ݧC�>-x5����n���,��XQ,�����Od:/z�γ��Z���Ol[��k�c�,.&�� �U��"���mކW�L�x0
�����w���MZ��P�0��-R) U2o�Ng�����dt40�R�r<�:��qݦ��L�,%]�+�ä��SvxA�mc��}��O�C�Φ�U�$�b>3�\t4 (gn���'`{�'7|�K��h
`h�F��[Q$*��4����@����d���55�y���=��$��n��NmgD�85f����!oc���_ز� 9L��)�)��1��G������ڈ�x�N��m�0e��/�-Ħ��T1ɝ˟p^"���� ²hHF.>M�<�n��C�#�d��YT������sۅSV�Zx�������fwD�ԼX�n������4z9���|�����e�2�hC�~L��c��Z�¢}�Ο�7o%�ð绡�p��}�v�=3�M���� v3o@�R��:�i�'^"������e)��u�����_�J2��R�d8��'�s:*�U[kj���_h>��gr����͛<K�>sN1	H�=0Y�r���{����$�^e`�E��"d4,�S	?��� x>{�_;�˚ě��������X�J��T2A�@�'�K�P$��Y���e�R�l�MR�$R�㺪B= ���o��EZ��8K��`�$�40���Cˊ@1\�Y�ӿ���'��-��e�Y{����Cv�:�m�V��o����mj��Ԑh>qz�'!j(�KO����gn4��JyC3�M��?��"��`��M}\����{�\{t\S.j�3Sst�߫��/�8T���3G����6�gj6����O�0�=�EЏP�A�v�#I�����>�����e�|��}�N	��¿���#��+ ��RY������/��W���K��\,����u�>�u�mUx�N��&�n���K�*ޙ{�L�e]]�˹���M���Jюt�+��^<y_e�<�[2{�8����@��AbZ�k٠<�:��V\����A������/�5EGg1c}	��=���%��~�ߍR��p�f/i~"�T�>�O��:�� tw��f�A/9�۽�d3K�X����mh
���_aߒ���;��^��˻1$~ZJ���}�rz�=p�e��w��/q��)�G��ބ��[�u��](�l��g��w^�8���tA��I
je���R,.t#�o�b+��ڔ�7����u��H<�I'�g�����(��Z~Nv�5��h]�1F�R�Ç�pw�$sC�6$K��q������t�ܭ��:Uq�-�AQ����?Ni5E��|�o�ڭ�5 �Ǩɿ睳���3ﵠ��� �ݓ��Aj�s�>��t�v;��\�����;�d��J֮�����P�8�-�{���Yz�OMGi��Z�������O�'�{�Ute�P@b��fO�C̷y�8c@���:�������M�G�X���6dտk\E�j����l�dʛʴ�/e@��0����o��8N��
���]x�)���5���!p~�i����-3���Р/8�r����>}m�#�4�1��A܍	;�0�-�M��a���%�� G�<����6��`ȏ5مt��u�WtF��{vhb�Ѝ10�h��	��A0� F,����4r�@;�Z��"ŎI�]�[e6�ޟ.�.�v�v����x}R<�_�)2���Ǒ~���ms!"�(>p��:g;������(��E�n*�����c�ͽ�k�mD���3Z��&��s^���p�e��d^�36,�sl[��S�8��U�+��_����EC������?r�٫�3�Lf��,m41��[��@��a��偳�/T�N���H0�F��v�6��8_�)"c�J+H�ǋ�;�u��@XƣF���������������i��$�ͧ.�<E��FbH��Y�t#�I��C����XJ�Ya�a60��p�:��޾�B���Ft�G�\��~_q��4�~�_Y�rt�/�D�8$��Y&d(�e��)z�po�sqA���/w"���/,�ܝrWC[X|8�����9p�LT�������O��7_�8��vd7�����~zN��+���E!�V�F��_���r��m�m{_&�z����˄�F�7;��+t��i��K��
�>`Xei^K������'N�Yh�W�D�&"��ٌ��yQ4%� �G$�K�?�yw}G9h	d1e�����-�<�:n0�x�;?���@������\ڶ�~B���l7���[A��ޫ'��g��љU~�B��㭊Ac~x����z���,ɼ	D�%m��廓��j"�x;X��|��4������]q�{fY'��;�,h��fe{�[��(!����L�b�=EϬ��δȏ��۫G@�Ԙ4�KJ=�9n<ߵ���hu\��uG;�d�/]�-�)W��NqB�E����d�]Ha#�?J��c�F��zZ ?�]���c,���VL"zlO�1*�&~mMݫK9Qw����S�K뎿�_I~r�g�c���m��)z��D�6֝������M�b�0���.�q�5�ܑ_��O5�>𩫅�'o"kE�]�q|�u׾����s��"3Wz���Dv�#N��G&qz/څ�U���P -+�k#���7=���Omݚ���%X�m̭��`�f[��̋�X�#|�!�������j�H:�j� ���$��9���2����l�8�#{VQ���$����I�Id:ȊI�.��)�����?����d30Naպ� �C�
���;:p,��׫�$`�13������SL��׈�j��[�Ƶ���wz���y/~X,�2v%Ae�[s�=�Bs�ܦQ�7�f�v�w�
���p=ח�N$b��+`ǹ��B2�;�،�ƛᲱ2S⋢����S�[�%���T�d����0�װo����>��}�b�w�t���4��F��kw��@�Ad�}�<��cmΖ�seʈ��O�w�\ľn����%eR��KLli� �5�C0	k5L�����I� �����A��i,茽YS|<�,L����e�hX��Tx�.�Rqd:��ғ��t��4�E����K
���ʀ���
b����AF.v��FV� ��Ewz}j�i��T�sz2Q��,c�QEY�e������lG�E}%���Oz� ��!���$_C���Q���ǃ�O��r?����1��6��W����u؇��L�����;u��zco69\h=���1)��}}�!�\׺m�28s�fVes����RNb+��>R����U�ǉ��'�4~ :*	*ޚ�+gϥ���S~v�$��-�Z?��O^�{�,��B]��@JC�����(�:�ެ�/V4-~�`I��9��c��
���ײ����X�k@� �m��q{&]�
�����Lp��_�KJ8�9�)tc�Ke�ےϔkl� �w&���d�UZ��I|��)H0Q��A��Zry>���ˊ˽�y1H���|�T�g�<����[�Xe�>mC���~�~ؕ��sz�������E+56Џ#\���L�X�>��d���o���/����E@Q��Wid�-� qt�n�y��+����X.mԚ��yҲ�d��l��B���]S"�&? }�䑑�M�޵�^��ؖwU�e,���h>b�?\�!���Ҍ��e���N1mqz^b�J��.��+D'j��(����n�(�O�[��;W�}����r��А�+����U��xI����������Q��9��[_�[�x����RUi���./��^��N��1=��~��;(݅Y�:Etl���(���� �̠1 �|$<80$K]j�ݰ6|`��x��L�)	o�td�<��P�{5OA�g��ݜ��72�,>�H�2Gz�x��k�2C+�/7�`��|�^p�fvڕ�l�3bVr���<]m�ø�W� ~GNV��z�#���"��LΜZ����1&gI��O���L~�j[��c.�e?�
��kMS��G�)�<e6နO�V�W���C�D��qL��E���ic��䯗����{�n>������˕H?�
��	�/�	�̽���3�i���:8{<��B[m9���=&YI�,�B��iz��<�=	���X�l����� �	�f8��1Dߔ�zޥ8M��T͔��tߤ������Kk�o��i��䳸���r���l?`� �5|��G�y#���*�i>ɒ�?}�'�N���2���֙���I����γ�兛dmB���ӟ�c��f-�<����'�[d�fzX��|B�����ϙw5�@v�c�~u�z�c��L�F�~�rd2\���d}��"�����9:}�I/w���)���L� �0@5c���z�.yϟ�c3od�N嫮��u�d=d6�囗��a�v����!�w�ܞ�)1s�u1�2�Ѥ��@�id�T�6�%i�Ef���ﴞ�U_d�k.��>Q$rz���gؽ��S�SQ���u��>��.6��1WvsKnsK9!��dZ�_��/e��$�wC�|��
�(��y�f�e9ܲ.:��l[�V��~�㸄V�IH�vvn��[~�/S���jyСl �jf��y�2>(�=�����&H\��%���{��t��	=�8��G֝�WP0?����/ ���o����d����ߋ9��\:��7�c�H^6x@�!;[?���v|�RC��1��R�& k�S�ud/�'3m����($U�L�'�Yh�����lCx�xƛ�֐���Q&\��U��TG�!-�5i���X��O��o<�B�u-�%�O:�C(�S��v�"{���͗���B݃W��W�)��?{���!��u5���>��7��dG]�r)b!+�AQ��>3q��VO����2!cPϕFv2�즪Ө(p���ӂ;v��/���S+�����J��?�0�Qj�u��xF�Q�R�c����HA:|�u�J�u����'Qe��7Ue�;"D�nL�f~4�M�5�1��l���2CX0��ݰb����E_�l��9��L��A˰��k�� �Ar����uzG�ӳ5��aQ 2��/t�j��5p�LF�i��YD�;�N
 �5chŏ�x>G'�hQ�9�L��uK�u���&���Y�t��[�f,J�M|�X��S�)9�;߄ĦD���C�Ԡ����a��y[�%��v���*�p)W�D�f�Q���a.XM4ף���{D�O@"V���Q;���������}��^��ɪO��hf)�gG��_��Nۋ�%��+��Tq�;?�c��'.��т~-��W��T�05)OpYփt�
L^��\�\mw�@���'k�Y���8�߄�Ғpy��A�R��*G�|M�h`�,�l5<����	�	h��/�Kr��"��A'�W������x���$N^,��0���؝�i����Xr�w=���*���Or[s��{�>;tI���E0��?�7��9j�R�p�)O=�f�U^�B&,��D°]w���O�tz�/�AoE�=<��d�%������+�Zд4����~�Q;I��
"�DM,�����أf������p�U�+�/\�L�^q���eGY���N��/qh�cKHwmC2%']�L�:0�Fe��f9��	 �&t���0o	�����)tZ�4�K�]�<���K�t���	c���߬�3F��K�(�<��%�bՖ�#J�齷%�@*���>�� ��#$�􆼝��&%���1���)&i��Z��`+w5��:ݍ���*f��ѿ�d�|?3,Ji�b���<^T����p�ņk��0�|����ۡ��܋S�W�>}>�y��+���v�#Ba�h�0��,�0�q��)�[�l���Dis$�)$>��7|�o*�X���?|9Gf?W]�ovmmJ��'ZW�HJ�bC�xٶ��\ \cNU<t�L���Z:ª���+��6k���v	�j�[����� K*5�`���	h�U7��S��]���1�o /���6kf��U9�J�;��Ӣ� o��`�>���4Ma�hd�`�_���2���\�Z�����ϸ���*^�]?lӎ��$�-�h��R�u�H�r����� ������bv�?�WU-�nV���d���w�T5�\JH���]XL徂����('��5ֈ�z���jjK�Y����Cr�����V1�rE����|)mR��4�m!	W����j{Z Bui(5w��lg���5뺂V~����8���k����#�ꜻUGe�U ��=}���+�U��q�`l��)��k���r�g4�ŕ��M��N�����5�E�1-�	%H0���'��Ƴ�A�{�9�C�����nf�,���cm2U��yI���c
.�T������7��F��R��3�u˪�d�h��ڋ�υ%Ju��}$S���D�	�&���,286X�5#G�q�>4)?{Q��.�ۋЎ8
�	>����:�] �̬�q�owZ�:�u��-�m݈8��� ������D�ñ��Ñz]i��l�"�[��?������k$��S׾���:�k"�
��w����& 	"T��
��۔�$T�h4/15�Z�Q���Fl�K��!An��ݷP~6���TPp�E9�W[ـVT�F��'|(��n��3ռL�e��}��짢�Ds��SK&��m��(�	t�j:ۦ"��.�m��aU�x�d�\��^.�����_�w�ӓ�dS�g/Cj`���_LB�:�m�F3�pd�M�C�����i��o>�Db��J��d�+B4N
��]&�;�ߠ�1C������z��.���l*3\���'8h�Ǒ)A���l)T��E0mT�᳑���;e���5:����N껫Wo�Yr}�����s9\6�>dj�T�xfd��^�=9��;��[��x��ONQ���E�3i�k�x�9�l���[e��O�4hl�e�_�QST�҄�����+�"�2n�j�F᎑�$��T��j���e�Q�"�H��wl����~so ���+����4׏�:���ʦ+�缬2k� d�M Bm�,�ΦMq��a��W��}B���BkM�;����;x��B_�㻢�>u��D�7�������ז�`Rk�H-)R��y�#N��	;sUFt�ө�6�$��Ƙ(X�葚�@����[����Y$m��Z�oK9?^�lgdOk� ǂ�
7?2StF4�[���n�pv����Ҷa�с�y�q#R+�)6�t+k>x�ѧ��ϰ�zQ���h8�55�sf1Qvk�v8�K�D�%�%!�.�G���|�HO,'����o��k�1��Ntdj�c�2@QY��S���^d��5�AH���a)W:/3�������P����=D����PK�G��CF��J�yk.��f��a�N�>�<H��(�z��8�!��M��vD���4Ř�Q6��Ӹ�	 (ԏ�Ea���������s	��"Ζ����!9N�q���)@���T����l]��i�;����u׹�K����ƺ]�>��7���e��^6�,ҷm]{
w��(�[���J2`���A>,����-%Rd}��.�G����QSP�R\�Ʀ}��E���y�)��)�ζ����֩����D~vO�[G�m7���<���a���H1���������q��������佌0�rdP�`m����c�e�O-����b��:�x�o]��C��ĻDs�$\Z+T��ij��;J=#F(����+%�(Mtej����o�U���e���"�%6q�C�F��q�L�__ѳ�y,[�o C~b�O��b��q��5̤��B���1:ZU�����|Ij�1&��xlj樝f��y\k��Ñ$�ʄ$��XQA}���گh��3��_����D��!h{h�zYO��l_����9P��m\�R0�F�y@�.!_.�k=]j��>8%�%�,]Ğ� ���+/Σ���̜�5����r��uL��r ��7Sc��:��0~T�p,L4�r�еSW�b�S�=#���Mô-��D�}�eؽy{@in����F������|��W��@TG�j�ͭ�9}܉���q�<�8����`�?X~-�q��U����%�D�39+�x��Rb��-^�:>�������;
"PყK!˻ER�5M)�r���l<�YD��w����p݁OZ).��A���S��s�D�Ɋ��ЁK!�␍*O-���s�{Ƚ����w�s0�s�kB�!&pfh����I'A%�1Z2�Or�\�]��j4�j�������-y%�%�o�K�b�H�}7\,��7����̡�M*F8������>�fM	y3]��'�zry9ǎ��sP���ђ�#�<��A���J�N��'Th����Wna������s���jѽ������9�))����l6�/!�m2D�mM��f�%F�d�#�O��ZoE�WQ;q\BP���u�t���)����l�z�7�ެ�)/-�s� �^�hH �����6�h�W�\Tյ~HS6��Y�ktl)��1l�z�������I�E�h~�5���殜;�;����i�衴3;�r�`υa�1 ��R���$A�[�%e}�fMQ)՝���hǉ۽��t��B���[�t�x/��
�����u�y��d� XU�n���H��S_,>jۥ|�?>@/������խg`�F�8�dy�2���_�bd��Q*2�xn:ۢ�d:���|�ޥ��L|��R1C9���9���;B}�l-.0�y������q�/d#�ц���4��o0���Tr��'B�����~2Nt�=1�[�a�Ù�bCx�[,>�M�lٱA67���,���oxĞ/����Db}��}�;����,}=u�_Q<`��|h���?����^r�3'���'����W��d#��o��
�}�`�,5D#��`�u����2�)9��SͧW��*���sJ�!�0sɈ���#Պ�1<6�]�
�I�p��0-EJ>kF=�f�;}��EaZK�����׀f�ʞ�8�_���'�hY��c.Ð��8�w���6~XUg��}(�I��#����r����c�fvM�Ͱi,�S��l�PH��������ټ�,�X�3|��D$��8��7��T�-��yBb�/"C�?�W�+f��T	�����T�0˻�^�1]S����`�Uf���l��a�w��+M�>!�g�e_nG���B*��H�G���d�>��/muZ�/�K��/
�̒�b O�y�[��,W�rkX��uT�B���S�.t�ĭ�3^5ݟB��@��J� S ���UM��7W������6�;aT?~@l8U�odK|�����! M/]�����^��u�~V��M�Gp%���}�����|�(�GTsJ��٩-�nV#����Ա����	�*�E�]Fng��"Œ�p�⮌Z0�C�V�qAj�Z|8d��viRSf�+;�r�������a�8i%��i)�qf&��H t�P����TL�$j��m�ޜ��w��Hf|Q46�V�f!5(뼕��c'nl�V���$^�`�^'�]���ۖ�X?'�W�E���q�[���-EtV�q	����J�H��/b�,v�p����3��=�!����hi�VU�4Ŵ��A��۹\��ɲ�F�E �+��06�C��#�H�1���up��p��L��|FaM�}�+�S�����,5Z�������="��ň�"��~K1[��9j�c䠥���i�Q�a��<_�7ft�8,�|�5~��њ���g�h�F>YvI���ѡ�왅�&����#�	�1j����J�xn��������-�=��J����=A�P�;�p�u)e�5Z�[�`���@�Ծ?��H��/��Fg�}��.�MM����{��?d����&�D;AF���o���^j_���e�$��Bs�띩
SA* /�e9b�J�P�����ԚY��iT�]n����|ᥦ$�d���?.�4\��M�PsE�
��E�(Q6���aE,�������u����`yd�
���e��7
�c�`��>a@x9$*L��_��w"��i�sؓ�஫�@�]��+�p�|A��'���Ռ�8aHfX`���|�H�W��/��n.{&cX��]�X�`�N\k��vB(K�D��I�ģ�n�"�zeͭ�A͖E�k9�We��d\���7�%uh`�dp`�}����k���Ԅ�X��/�U��~0�m�z�E���'��Lϛi.�O��S��t�w��J[=;ks#pSi1�����Q[�^! $8��������+�/*��ʼ�Vu��H��U�F�gK��軠5���5,]����}T:���+��%_���;��-�n~_���WO����^���j�1&R�G��#�.W	 W�YdQ��)�[�c��&��B��|M��*RO ���1��#��y��l�j�e;Y����%v�@������w��!�	�hc���d9�+m�-�TW�x�zkR���E΢j�5(U�5�|i�DOy³q��6�QID�v�6꒿�h��!�M�T�,���l����*��sd��_��X�bJ�ٝ�)�vQ���`cf�M�}���Q�/�d8�+)�/]���hfi�zox�Ϥ�c,ą�]L�`A��&���|��5i+m�_��o���א�qZ�������J�����>w�I6��ؐ
1t�=O�l���������ۀ��Q��3IJ#�ӽ��\k�b����rRϲF����fλviȌp��gt���I�.E���!^���"�zt
�����g�w��@G��v#6q�V>������Iߍ{^��Δ�<����h��yŠM!������(Q��E}("�z�����L��q�lJ��'"�v0"G���gm�+�pC���;�jTx��G�N���}l�Y��w��2�0�;��RF�����;f6�S�G|����ٗ
��^�� ?y�̈<&����r��y���e2�U$���U_���4�*�
,xH ')_��N-� dՀ^��vg�����!]���=66K���]���A��n|�9т�R��	=p�8'Ѳޫt��W��jp��u�d*g�Qh�M��*d��42�n����쓌���
-��ܿ4�>
�"OIȆujp��/�+���@�eJ$?.����u�n��J?P����z�͚΋�ss�o���T���ٞ���k�����ބH|���4Þ�h�,�#��ynL�q��A�`E�A䛵ܪDUשZ�8#Y�z��O9��+d�N}3:�R�p�|y�O��G[۶�����<�B^>:��dxБ3�����HW���S�<|�^���<�-F]�SϨm������"Co9�����]���g�'!C����X�����o��=�AQ&^A���8�ޥ��}�pN{��Vo�� r��@I�c!���br��䬛K�6�H�cb@�NS>�?cոx}}�уh�]Z�vGk����^�)lk6w���!�5��2Ic�99w�u�@rU+�g)�< � ����fGu$dH��_#�Մ[��OP	��`�g$���?�Na�r�ƿ	of_d�bVu �M�:�lK�aKbMy��V��0U$ ��f]�¢ϡ��p�@���6!�V�>/1 
O!;u����?�vV�A�P��']pz+th	��5o��B��l�P�ސ��58{�=醻[1��(}���!l�@����cY�3k�	Q*�KK?��1�d�&`�g���F8���)��?���KP1� {��MR2���bIz���/�"+�ُY�����^�M�[Fo�{�AQ6�(�oi���e��B?��o>I���*)��.H��aΑ{(�=$BP�8**
����޹�ɖ!ݯ5��@�9�>}���}��,�X�y#��.qz�̧�OE���jI^��}?���x�Jb�Q���@�Q��Ĥy����Luj��?����NG����\��r�$1E���"�O"4:�>���'�q���k��C��z*�l�2S�����>*Sǐ�i��-]o/��$NE3ػ��7Ф�+5��2l�x�jy��EF��4�;܂D~�vf�W���呺K�ٚ!P	���H�A��U}į��G0�K*=��}k���$�x��V�y�KN���=�)�����X���%�5���;f�c�o����J����¿��z�N�����k�g9H�!��R�/��KqU]�3b��w&��Z����Р���X��d˿���s��Qo8.h�9�o�֩��"�!�}����k�v5��1d|ωEW�W����E�	q�!����l�ŀ�=�_��u�%�":��dh�������B%������Ym��>�/I�̀n�ݔ���4i	���+0����D�'*@�����%���gL,m��8��
����d�����t�f����į�cüe��	U;�إۀǲ~A���v
Kjդ��ɕF�G�F7f�ҏ�	a9D&��W��͑��@�O��+.5N#-����n᡼#�gQι��;iR&����9+���*#00y[~7�����<�)^��k�ޮ������d	W#�Ҭ���*�>�\�n h5}����i��m�|���Aؠ?�F�G��� ;���8ݲn���-˥����,U�,��w�����dj9���aai�P�N�&��2MC�������,E�����NxlA��HH�>�5[[)pz��)����w��m���g�4���&���%����eŞ��g&-t��6���������"�P���Ba|�D�'7N*0Ա���/��}���"�:r�Zo����^�a�
�@�E.]���ہ�ޏ g�}��^�M�O�����˹k���8fi�ܲ�O�5kY
�э�/�Y��F?<;(�դs�!�J����'�/q�:c-�>�:[?i�6i˯v�8t>�'��gs���Dn� �&��s��ڐY�k�|	����5�I��9�ɶ.;��,Ňo�S:�5-�뗹8].�goO��,�����^�<�ey��ړ����~�]���eYh�t��n���hj���/_��ez�9!��s7�A3�μ��{\���4��g�7R�xU��6k��\��V _���,�4SP���`�yȒ�b�\T:�K�W<�nI�IHD�3Y~r����ca힋�}(����TV������t
���~�P�P}�u���oa�W�O�ϰ t�<|�����5%?�5������%���}�M�k=�P�����m�+2��������i"�^�./V�'���؛���o��;�_��4�H������f����:�1�["�k1��X�{�s]_
�e�ۧ;AL'm.�$LN�I�[Am.QBK,i���mwҬՐ}��9�����M^��ꓜ�(t���}l�3 D�A���� �i�Ub��j�����}������ĝ��-c ����p�N�D�<����3<Zj:~���sϏ��?���E6Ndڎf��N��x)OK��4����7�k�o,�f�ŇG��"�ӿ��$w��	u��0.���}�Ԁ�q�����F��'�N��@Eb:+���](�������+�h�o
Y��Y��9���is�h�5|������k��NtR���ᡫ���^p�ʖ�*g���r` Ï��l��Td�ڈ� �` ڳWI����9
�(e������_�%��β�i_�����l���ƙn)#���`���
�|�#�!Ig�5���N�e��ޘ��qM�N�p�=$F���_j��2o_�M�/p���y�SFi�wԈ���u�q�c�ј�A�p;ӀR�S2pl�+L%@�:��.f�l#�����鮀�( ��iC�-��}��B5S������1%�ʲ�[�t1�`}|��q�WI��Y-3n�oI�hڿG�m��$R�kʪF������>?;�w�����sx*���%�(�u'��I%���S�R_�B*����{��4O�%ݘFmo-K��?�&���?���\-��-j���;�)��q)2E
RPh$:���:�Az���>���M4]��#�3(!֛�a���L�ՔH�V/�lu��y��bn�1�l��sS��\|��ac�{����\��c��1�RΆSU�uS�_��8蓎��r�)�A~�.�{��<�tn�}8�M*v>�T���P��<D%��s���](�:��̍�W�궰'D��ʢ���v{��SGT�#��Sm�EC�p�2 ���|.�B�w�(��Բ�)Sa�툩1R�/j�kQ��NF5Q h-#.N���� ��UE�U/��Kc�A7N�Ys'�
Ǖ����>�A�?�C�J��(DpL}��uʭ�t�;C�=6f1ss���$r\���wZW���(裒C|!���zm�I��v�F��y�dK5a�tiC�� ��Y�ﻹ�	;�rj�#�2[Jf�a�#$�ȧC&z�����o%hొsq0�{��/T��'.���~D������J�A<��a���?}��{�������<쉂�Ee�`y�*��-�e[9�b/M���߼۩n
}\��a%��OD�借V-{Euh�.UI��
� �6�R�<9w������H8c�,f����ɡg�3âUS-'�ZhpD��N��b~��!|��'�UZ��b��NQ�*�Cs���ΰ&B�*�ks, ��%oo6����a��M�ڣ��r��qc'�lgCRT��K�Ñ�v�"��?��S�d��X
 0?=����%J�#�g��a�y���'�!4򌋏w�uK�#^w����?fVFl+�,��H�J�^��.;G\ۂ�~�n�%y��@�y+>K2��{�ZX��m��`:�[1����樦�V��S)��w�����t]?�G^l����~�NS��S��sM�a$G���F��푢�pF}`M���t�[�Nٱ��k�Ț?b���BK"_a���ڡ�����|�s#i`�&.no
�~�4� j��"]_.zI�]`}��|���2���a~�h]�z�A���c��W��8�	ׯ$��T�F&���L�� ��V(�q�Q��Ӡ�`�?�&���f	��(^_d/lXe$�~���#q��>�h-Rd�ޠ�Q�R��<��5A����NYc�Gx)���V�O@���A�w1T�Ǟ*����.������߱�i_?�-3T��PD_�NU�������V������AfL��H�v���Xib�5 ���h,fۣo3"��bzFz^Ѡm�`9�	�"��Zؖ:{-�o��������G��&�BU�TƱ��ܷ͠}Õ�������d:��/�*�\neW���eL^�ĭmh�Jq��/�s{D�Hiz��v*<A��_W%v �A���ϐ�B3�j&D���;V�y��7�A���)�?P���/��|NtX��6u����
6l#���(�:��g��qX���ͯ�T�]�5�d��ύAQ�\� �Z4,sm��=��Ab7��R��j%�1�J���/�1���mAX��z��k?���t�F%_�'6�W��8�"��w���O9���ޞ�e�v{�����au^*͢���&��f�K���?1ahs�����렠ka[v������GJ��������2["S�/S����ݫJ�[L�����d��T]�ȭ�WU�0j���0�f�Z�'�H�lnņ\�����V^/1y�U�r�� [�%K'A��C,<�伥4�ew�c�U�k��A�7q��Z��䯷���T�c�V�y�
��.�;�h��#�P�J��I�4�z�܁�� ����qQ}���0�t#!ݠ�t���H#�Hw��4�]�4Jw�4 � �����}��f�ٱֳ�z����l�[{p���lek�!�_8����ym���Bq���,�"��vr�M�Q�|�U���Od�h\ҧ��Ӣ�̳7�*5�;dP����:�v׹�|od�|n�ž�e$�~�"�1�qw���H��>��j�#��J�s�E'��~T%}H/���56�/�=��2�����wL�_'}墄��C�F�ۨ�I�@���[�w��q��Nb���[��麱s���H�z���p��/{��&��P�09��Nx?[���J�6�� )�$O��#K=�M�C3P�r/�n��:�ov7��cc�n��CD��u��v�0�^>)��gm�&Ŧ�=��0�/��u���4�7���^����#����!�6U�،"k�DC5�8�8����I�s����^ƀ��-ػ�7V�zfxt�}#S����r�����=���ů�DSz�D.ũB]T���Z|Ư����Q����^R*��ׯ������������(��ӎ�3���\ˠ�r��MK����2�N��Z��>>�c����߆���l��~3 ��p%֩k�o*�s89���&��A
�̆6&E��f�s8���F�J<gvҫ20���;|u�Ə�����k[�$��8[�u��'��:܎���З�Tpq�o)��}'B��u4�8**}�#��b�����u)�����a�bG��u�t��Ѱ���B�7��mS~>�B�+��g���@:��j��f��=���ɋ�'���>_N|b|�Q�f6�V�R���9T������g�8u�f��u�t��o����'O�j�s,��q����jvJ��%���O�{?4M���W�k������n��f�Ƞ��}:�o*�?�b&s�)��0)�/����� �}�o���H,�o�Mi��Gj*(C����u#�|���qGQ��rb��E��:;��۟�'�juY���)��h�������'eN?�gw1L��-LE���E�ZVð�%����A�8K��1����b!%S3��+Q�ݔ ��:�ηmd�7��"l-���ty4���������Js�B��Sx��abj���djQ,��F�Ij���f�$Ks��P��~K��_�`�F��>wI4�����x��|���Xϛ�@�]}Ru%p�e0STTo��pC[�5���׫B+~������eyK�vrC��n��B���L7�m�z�E�[)�WAx~rQ8�b ӿ���}pHb�ѽ����(~���o�#?s�s�_����X4��8�x�A�3SS'(��(`{(��y$D��o�\������]Д�t�#k���+�Le!�}����V=������J52�J�p���"Ou�w�~�S�W�q&'K�(�܂����j
{u:q��+ݪ���?��f�=R�tN�b&%��<;�������쩮䣇�/i�|�٠Y�`,BV�S�\��4/����@�J�o�7&vr`�m_�[Tebϣ�#㊜�����B��Zm(���p�)c���P�L1"����o���4��{�c8��N舀���&��h�4��T��������
]ϳ�{?�H_-50����">��.��&�U�%���� V�.�A1������F��.8 �W�f+�� !�u��j��^�R���eښ1�CB��zDf�}�F�7����}�_#�h����(�?���,��u�W�)���?Û�i��ȁ�%��B����{X�
Y�kʝ����M	�*_�I�g"'C�WWX�
%H5���i�D��PɳP��dfs=[�v#�Q���V Gn�u$�ß�@�I@V߁� �B��t�C�V@�n��xN4�j�}�w��o�;�K� 쌖����L�uqr�^6}�sqX���u�C�8s⿴������Ž���d��N��}�V�v/0��]Q��!fX�8TB��y5	]��ytl]m���L$˳��_���v7}��A1\�MX��Np�SNNƹ]&�>Q�|�@i����L�cZ�qSTY4)�Q4��3|�5��ϛ���}�'����r�l��o��\���ڻ�ϡ�	젳WFS~�\a�Ls�#�q�ab.��DcVAe<�q��-��%I���,Y�z(��m΍<�wC��~v�˃ H���|�a�b��,�����|�D���"��=	g����_1�z�����ag�k�X�cI�q�w�����w���e2Ɵ��CP�.Pܗ���R:�:�] ػ��9g��lh�^���uݞ�����xξ�Yld*��5�$Y���%Q�p�����G����־� �%0Yy����P���_��#��d7��!e�["��<6/�����Q��A���~Z<��V�2,&��d���!�����}E���'���s̢EN���Ƥ���t �D\؈�n�8y���"d���>[�l��2TJ����T�c7����_��=�d���Ol����z\t�g�e�]�R�� F�E�{E����GZ�w�����*�%�qˌ��9�T}����9^������aR6᫠�Px�3|ZW�]¼�d��6���lзtx����[]��2�G��q���w�
���}�8��8M�	�:��Cs(Z�����J���������\�=͟�m��.�$(���|9�Y�8��yv"��$m��H�w�Tn��E~y�~�5w��~cGC�<.[k>�ٻhh��~D�h��'����T���K7�Wj3]~]��9���hr�W�D�kc�=|K#x:��S��N����,�Ԣ)����Z]��T�6�b�XҮz~�S��z�_�z0�P<�"ˍu���t��q�+T��HϾX�77+�ǿ����M�8��s��p���_]�=x����!j_��rr��/�fq�s�"MՋ8��:�A� 1���#��jƼBA.aj>���p�[;?�����B�y��
Yc|o�oWv��JH�	�����p@�*�����?�}p��?F�N��?U	 ģ
���13�w(�7�\�|�{I\}o��s�a��{?��9ϲTW�
:`{�d����b[�f�"�NN�{2���t�'5������;8�^�����iT�8�O����b����;����Yׯ;�9%�Xy�̫�GY�wa�����O�Tg�q������X�t����{�!X3�N����yyעZ^�Q���9H��R�ٍof64�
�&�T�ä�}N�q.���o�t��E�P��j˓a����n��6]:����yN|�f5�z���[u��[*�F�c��"����Otǳ�g�8��gOi݀W|���
�������:�<���&4����X��EV��!c��������R-�V��U����������e���1g.q����N�S;�uRW�nu����E�Tz�R�+�7Xܴ�����'���L�(xE�n��&���3�C/inGJ�A�����(��P�RGGez�~�60^ͭ��Q�[t.ѭ�b����Y�!�8B��r����	h:*���q݅�v��*�*Ǐ�)���j|��Fyu�9𯚼XDt<��ф�+���}�%��񚚍"��Η���;i����a"�i��O���ʹ�w���*��H�1~�ڬ�[Q���,�`l`s��"P<"ݲ�'�Uϲ�����FPβ�d��[���Λ1��Ie��^�O��o���]��/m�Rn� C� �����i��d�&���K��`,!��۝~ߕ���_x�7�D�s��Z�\�>�?��mj6]���贍|���ﺁ�̣�`����^p��{��q��s�IX�c�����!�ѿ#�˵�n��L���m�l�������j�ύ�K��� }���?w�f�(���� U�������F��IՇo;>z�/�jG
��eW�"�(�ē�+Ƿq�1�+,��-��{�v	��Ff��C����a��U�p��P���O3�2V	]���"��F�~Ss��?�x�?����䒛;�6��.L��ݡ1�f�*���*膾���oL}X�28PK�s���0?o�+�`�������d�K��XY������Cz!��8�������A<�nX���@=����*�kab�N=FW���3| Ō}�h�
]Y���>ɸ_?���S������b����V������Y��&x�˼���ۭ��u��ȏ �������Q��Ǭ�a�W��Bg7���s!�3��I�W�c�kc�8�+�Te<h�R�BcU��yd�Rfc}�c�$T�DK�4���l0i��g$�<]ot�G��*�.O}�x~�z5zo9D`�Ġ`�Y�5z���Vt��YԡÄn��Ir�M��1���t�����tZܮ�*���P
�������J�h����Uj���h�!��CL{�:^�C����gl���}��rSr9��N/N�i^HWc�RU�`�8T���龸��
PY���|T.d&7�a��.�΃oIÎ�3 �X4Pm�����>@�o7w�������$����,��.k?��`�Cl��AX�{�3�/l��ؤ��H��0���d-��xy��K����X<B/wް��7+ϧ!�sx/l�Y�L�����P���X'2���'���9�����JI��p�8��˻J��+D�pJ��A��Y=K2p�(��꠬�HX�I�#�[q��l�cܓ0@�?(D��E�П�����A��\Ā絥�����o���8�ź<߾O��c��}'���s�E��~V\�aɮ ��pd��7B���0E�P��O�;e!���'r@|�~����w�yQŏ�N��v4����I*h0>�4�
K?$�ȋ�Ր�eZ{�?$�;��9n2�(vDx�>����䭑f�s��t�`�Q�:Fq(������������d(���������	�cH��W����3)�X8_�7T�ܧ�,AIP� �:���j?a��� ���
`����S��I��"���)(����xe4��|����D$L�n��wn�Y%�����-|�i��\Ďވ�&�P<��`�[d~]{'�گ��1Y�"HY4xm��N�/h%ǁ�o/��.Y�㓲��,��L��Y���3G����Z�Z�2~0Alv��u�9�vlņ����`G8�G���zI6C�b�����{�K�?��Q�[qb��mz+�Ĭ)��?��aq/<�ä���X���I� �{g�h��z��Y�wD���V�w�g@��P})+�l�|a�l����� S��@p����uL�� �������"�뺁 �6��7�jN�K^c뀂W�f�Y��%Zl�2��R��jk��r����<��.I���*�-�Z�@y�d���I(�n{L�|d�8g%�[L����C܁�Ip�/T%Z���NM��2N8�K,�h<�W%��|u���I����â�E��;�/�,.�&�
L���S����t��.���@99q���̡��9�nIgN�Ӷ\�K�'h���kT:)�����#z���������?�g(����et���e[��O+�q����|�.d$�52A7�C�5�z�/�n10�����`���v[2�u�Gm�?W�uu\��E��"�+5��ÜBI�rK��~4���H*�)���J�W)E_نT��
�$�D��$�KF1���������m�))�xq 0~����ĭ���oC���z�* �>��(#i��i��,�~��.���p+��N��#���b2]�OL?�����ʍ�2����G�G_�o��]����mkB������m�%�4"�T[����u}-���YuR������9��
)഍}��[N�2�Mƀ�ˡ��~K�7lN|������7)Rh���Z��d�Ϟ�69cX��'+�)::8���'��y�We��*�������핀�j�Yν@�jYt5����Ǐ{*hG�f��EN:�Sn��ޗOQ}����;��;>1�#O[Ky�hR�G	�]�}T��d��v*�7G�y��z�BC�s�3!f�-�{)�xҏ�tL�@-��Q���bO�}n���.���~u��8������eaw�٧o�Y˾z�2\((����u���Q:*�4�4�y�ʴ�k@�ǲ��`:��q��R,�����I�n��ص������^�1��έ^�bd�
�I�2�~ms��Q�JYN!�Pe�ʋ��A?/>�;tT��S(?���t	5�����9	A�i⎫�(��Z��W�㠒�ā�Y&f��A�`�Ш�LM��P>/�j���qU�m�� �7E=ڭ�>�6C���i��2��=j՜�+�"d��vb�-�B�
i7�=���1�l@s�o>T�y*"e��Sr��!�wjf$%����O��Zu�#ֿu.G�Z�WYC|�|��%��C�����U
&�w���*��&Сe��tn��}�E��	��R:�-ɗ	*�yK���������'� �/Ǜr����L���#R
O�����e�˝��g�r����ٓ�T�W��'˕2����F�B3y#�ux&�M5(6q2��r����*���F�˂̡dn�d��3ˬ�6�� �����I�W�N�����0���M�h���5qr�M�:J�'���瓙�P�)�4{���=l�t1���&���Ԩ�H/�����/�]�,�������a5Gp�@�����j��zꢲf���G���� H�|H���ӛ�	�~2��5�ɺb�wn)��(��
#�륈�S.�6�>^��n���(u������kt+}��M���,>
����,(�{9��7�K�YW>����ײ�Z���):�)�W��q�5�L{�`Gw|F�X�E�<��yY���=�L"1����aR�m����a2J'�����Su�f�/a�=�c�-�q���{�� +7�_��.B5�7W��@]���G��ǡ@�O �ON�Ĥ����'����I�����9�V����C�Q�-�-� �������0�v
�Sֻ�q�����˪����J	��c�f�!�J�-N��`����v��I������&�1�'���
�M���{�{��]�o{Ȑ2� 
��N��E�Y��t$��x�N��<�A����M���/�ػ�L��>�ɑ!J�n:�--e�rm�3�O����C��y=H ���jdR�ϻM�9_���KMf�k��i���I3�V�p���r��p��D�ߡX�\Q4���kOYY�r࿝�bZ��F�lU�i�8����9;��.BU��[�$ w�42W�٪�&�+�s�J��#�X�������f�/��* �UC����Z,U�5>�1�w�n0^�O����[:*=M�5\h"m��J�e��++%��t���t1џ��d�\S�ȅ�
4�ԛ�`5Nb�G��LP5bw�������{	Ǜ Y�+���q��W>�ш�Ox��t���\�d&�.�ۦF�iab�dy.$��B&m#�*��q�b���3�2 Ќ��G7��AObȝ#(-X�3��hGt�UU=�n�r�ƀ�����_ޠ�ℨV>���v�ة�[J��)� �-�_˰7�q���F���L�2�r8��jd����3S#���	6�J)тC���?~����2���ڱ���W�ŕ�ߟ- �M�vQ�-�$�k"���dc���V�ˍP�q\7���a4g���ptk�8_KX��6_[�8e(1�/,ԙs�p�BB'�_��g��ǡ� ��c-��f	E�A�� �@q�t�&��6*f���vq�鏌�����lن���У3����{�A���
,�aG7�:�2�/|������Z��ZR9��C͋�����êO8�X�K<A���Fp������,�����5P��V+'���(O&�bNhP�d�6�@�o� �y6o�-��iD��"��{�-E��\r ���ع�FHe���O>|�טG2���s�D>_�u\�_��A�,^��n��ĵ!ff=���b����;ۮ� ��ۯ���P��Cž�WӮ�Jt�	�R[��e2�]�_����h�WU��6+B6}�<S):�m���J�2�?�>��A�ؙMp巣��D�)f��������&I�ר5}�h}Xnu����G��ߣ@.�(7x	�4���'��p�:t�_��q݀�4D�`ڕ�(����RW;d�̌�yX���hX�ZUP4����S��)ftY�4W�Q:��ר��z��"O٢��foo�����y̤c��
CW. �����!_
�+��j&����MΠo!ؖ%��Í;xE;�&3�>�Q�e�II���>Wi�Y\Q?��μcukS��es�wS���z-6��A�g/9�d��N8zd�~hٽ�xx��@���@�(�/��P* ���\���QWWd�(D���jХo���ػ��ms;�����A�����/�98t/�b3��Sy��E��jo� 05�AJ��l~���okuH������p*o�سﲜCc�1˹����ǿ#W3Ks	�"׳0ww�j9���&r�B���hݚ�D����Ԓ��C��"i{m���ˈsYlW��d�N4_�9��KqX,�x�49"B5����N_ʹE}�c�b� ~�#K��C�RU��w��
W!�x��p%=�9B<�a~��r�v0Z��29ۀ��ER����F����
�؃��4,���ߺ����kKx �ŧ�$H-@0ݎ��܈����=�����nFO�A���d���7\?j��y�
��8�̆��`�H��������M�@���m 0jd�@��	���� �����ueE|���ĝ@��!*C�H���'C���q�a󱽃l�V ��he�j�E��Y�*Gc)�.#�?X�O ����"J�R#�߶(�K���FT�/҉pOS�t#)K�T�����l�I'�WY7D��x�iC��M���>]!���P���z�1g��4y��!u2::࿍��<ko���`��l4��
I��d1�0Y�c�S��(�\�J���W@�@
3� ��'��^�k�PßX���X( 74����f��N'�ۍ5����L����:\LN�j��X�rYQ1>�^MJ��~�F/�֏P�L��kj��C2C��EA��m^5��q~���!����a����Z���ӕ��斥<SD-�f?�r�nZ�7��94]�B\:�2R��,k >3�!$T���@KX��3,���R��p�����0�m�:��fK��c�Y�����B��0�^��x#�!�!V�_��M7�|eQ}n�w;|5���kr�\�|�x��JAE�C�k	�C�:9d��Ԟ����I��x0�B �,���vÆ�sX?�Y�Y�v���O�f]����:=/l�x��:������;��V8E�S]�j6�W���y�̈�F,O���+�J���B��F����C������p�E�B]��$⢎K-�Bw�*j���I�YUJxK�����K�x�5����;���|�ߤ�M���ݜm?I��l��KԝCp�X��l���L�*@�����e�楎*�l���QPsl���_��;G2�'6C!�w�|i��շ�x؃��%6o~��MS|��m;�J(�D�H�!���B�m���W+�\�Tf��Amw��K�2��|�������"e�,VB���i=T�G�%�J	4b$���2���@�u�)�_�4��9t$�x��K�C�ZJ��+b��?w�pb����wI<-�*�	Ke�#;�U�]֡��	(0?2�a�i;W<j:�X���b�+�t���e(���i�GC`>�m�$z��<V�su���ܬ|�w�L �/|�>�6�&h�8:Ė��qP΃������1*���(�0cx��K$%���%s�N,��xHR0K���z��X@c%��O��LB:�%���(����f�>����Dbe-S��(y�?TN��!?� H��_��r�}$�Lg��B7��A�-�F�uW
���Ǩq�@;
̶�� G��j���W�&4s)r!�SiL��	a�M�U�k6C!�9�9�O�/#�ҫ1�Rś�{b_t����y�ʡ����C {�;?YTZ��Kc��!�	�/&�5�x��+���6�k' ��{���*B�Cr�ρw ����:C@4O����iI���yȎ�Js�"�c#�Ɏ��
��r˻����2�����M��_}�j�cP,�/�M�J�IH+�G\�\՗С�YF�R8_V@t���uE�O��eD<6��'x]+�d��,�&Yp�x+P�fN�̡��}�{�{����&$��,>�����ǋ(.C=J��|y�c�y�?�(��eu� W���4͑��	�<	9�����1i.����������_7t����uYZ�׋thG�}�&ȝ� i�RO�y,ܜ�����~��E��y�F�/,���K\�.�������Lڀ��A?VJ�W,P��ሴ���� Pk�T��uH�(&`���2h�cCH����w���(��N$�	F�������H"�n����2k�|=��u��j	�����fT^r����w_����%`�������P�WL�@m9f1��ͪ�G���m�u+��EE7�,�T0O�]�Z�v�`���i�~�|C )0b��!��0|�" �o�ʡN�R�,��aM�p:\�O�������p��\���$��q���1:�m3=_C��Vg�����  /9�'z=� �	�=_@
�0 $�]_�,*�6��eQX�K�^I��������dYol�:]�9��������8D��,~�G���3��S�ϊZ��q@|�0Q� ���}t���Q�����/m���r�uv%B�ri�>nB��� D�ģ�6ߢ�@N�o�s�f��MK]ث�#?��7*ʱ��y<���I�0��0��·�;�㆐�|� �����,��^@UC3U��4gn��K`�*��Y( ������y��x#1HtAUbAԔ�&�q�{m�8(<�{sH���5����a�ׯG	�D�e IUy�<�NP�q_�^���zZ
j��/�UV�[�٘L^,�윓)���3S�8>�Q���T|�0tEw�V>*nj
���iL�N}�2�ɿI�gL�����E4��	ȩ%,~�3(Z�bR��/��B;���X����\
c�͍�#��H/��?&��B���;�4.ĺא�`�,�s�!h���@���W�o����׾�c��Bѧ��F��C��Ƌ���ۼ�$K+uAo�}��įtA�#6;<!?������	���o�!���$�t�B�)w�'6��z��ɏ��R2`�UM�b,A0%�@������nҋ��>��Ht�r�NwԀh06q�:�r"�Y���)P��Yqk�\1����>��=�X����.D�����\v _��кɑݻ�]��
+�#.�pǛ�51S�u�S娴P"9%1��m����P'��&i� vv�Y�`C�R$ 'W.l,C���w,��hu�g�>��4RgpS��bu=�"�
�8[X��c�x+��ڸ��*Ǥ%fl�vK�* ��r_߉E�c�2����=��h���
��kni�'Y�'6�|/�&\x�����+��];i��}�|M䷧�aȑ�t�n\�=3��CX�.��� up��(<��:�@g���IigjP�ͳ�������ʟ`, ��	ts���8&��w.����K�a	ͬ����g��YGG�O$�p68����r��k���C�*=59��;��sL�c_c��e	��x8?/�����:[@��^�a�$ht��HS�cN�o�����#6�&�h'�\���?F�c#7a���}���n �{C��+���^�(�r�X ���h콻!��!���B6v󓞟��<svAy.���-Klդ���!��β�����O���p�{6{D>͗Υm��3�|���YAq��Ȣ�P�uD��i�Ħ^B�A��\��- �)�|�'Zl���uL����@���p�t8B�/n#�b��x�(M��r�YOd[��KS#��1���۳�i��ށ�-r,$%hw��Ԥ7!����F��Ua��G��~��S����!kEK-��!��B�-! ͆�X��RM�گT��l�; �h�`��ի��k�n��K�榧q�v*�ʰ��)S��W�W¥,�����ީ�|aw� q�sٰ��t� R<�e�V���yy�s��|P���5{
H?�����%V*�1-�U�JJi[��*M到�x��c�Θ�ʕ������|�x�'�S��o	�7���YM��s����kf��j� �H�]l�3��C��+�1�����j����������G-��}	L]��!���J�2��/"�6�KE|1W��ũ�G��"�-����%�3$V�G�.���-y��D	�y���CѦ7���xd4k �ۈ7t��w��
��+�G��(G-fi�/�f���@���H��G
� R2��h5��9 ��6P7P��Ѐo����m'~���W$$)�u��
�D�0vU�ý�9�yj�g�r�wO� )Eac�?�>�Xߑ��shf���
�K��J�u� �pM~f���j�'ɫB=rX�4�s"��u�|K�e�����k�S}�F$�+�����aE'f%e��y�'�S����4^<�\����t�|=��p�G�=q�"=���S�?զr"�E�IC�dq����9@�M�mUkO�ԹM뺕�B{���H�:�L��n�Ef���e�����_�5)	�F�d�?��C�gD,]��Ƕ6�tVw���[���6��������H�$�oX�r�qI`���ç.e�Ʋ挍-�w_9���;�^M�Lifa�/�i�#nRH�-����ѓ��A�[���J�^kC$�]�
=�7YWLUӘ�a��oe�b�\KE�h�l
��jV7��(gV~"n��Rn��W�H�ֶE
چ_2+)���Ij/��K���t���Y�\����Sg=���|�.���+�է.ٚZ�7k�0A/� -4�i�mV2,":_�������Ɗ��kf|�*qw1�y�:�r,��v��ݔ\��}�P����g)Hj�8y�6^�e�-f�9:��P�vR:����@����hQ �_ډ���4�Ц���Aj&ס?E�e�j"U�;џ����e^�`2��8�*b�Z˱�$V
���K[�C���!��>�ޤ �+7ܿ�Y!=�P1�:��{c`���ݭ�]}��[B5��H�v��ԇ�t_�D��@�lQJn��ŭ
��R�Z�����W�H���-���OVU�֡����BPU`d�|z����8(���0p!/��ͫ%��a�T��af�Ӹ���aW�����x
���ul	��l��&��z�7ӏ��*����k��%!Dk��|��b�v<o5��M���e%���}��|�&Q���>6��ئ���@zM���\�x�ݞ�9��(��,�ߦ��]e� wц^�D?o��c�v�Ґ��h�k"P/�7�v����������X��)�D��7��tm����U�˩�|Ǒg£�%V��T�}LT�xB Am��G�-�s�
t�:a!�$��N�Q5����c�$�c�a��'�3vx�_���͹e_�B&a���>�<߶ P;52+iL�ׅ�N�:�;�J�������%;��������ZNn�c=���3���i(�� ����� �E�{ns�K׿�Y(g=��3�|�X��;tK�ǡǪ��<ou1��ܟO"���][������l���G*X|��pZl����]���z��Xq�N�ٗ��%U�?ۨ��W(��ܨK�k�`~3��6�czI�f�?5�^�튮:�4�v��9`�h������{����C�d�g��+-�yB�\�N�`D-.�>�Q���D����TKKc�� d��H�Q��n��3�Tc��R�r��}���u��h��ݗ$�P���V���?�ڝ��w��ɭ�Y\��h����V}���������P��"�
<;pq�4�<�#s�G�~�U;xMqҁ����]޵X'��{�*�����5�f<&��ӳ�.�{D�ߕ-?��@�9���n�$<�<�4!(I$؄��XSS���<�	R��R��B����rX{×���9H��츊	�������{/��Gh�@M�T�cN�X|�@aߴ�����	��Z�{��L�?�0�O9�+{ɟ�Oph�)p	���h_�bj���2ϜȠyab���c�)S�L����+�SK��V�Ч����;������)��%�z���#��5_D�l{TWk�g�G�罉������e�.u�i)qKQ=h��3�.F�@c�Y�[t�O~J�R=���4\�=�~z�J�x���� �Ϊ!����֔�e+3o�˃�`��͍Q:��\�9�^��2 ҂j�vZ,h�(S�� :La**�>0�8�#�D�nn7SD���Ֆhq? ��,�&��,�����?A�W��,��K�i���km��n(�)�L��ğo�68�KP?��+�Lݨ#t�*�yv�d�3��d�oʫ��5�]���V|���(gbJ�!b����?�d�$��b�.�^�$�;��Moj���C���퓝 �pLr�r��%�3�6�L��� \��,�n5��h����]���>6�d#��%�>�3��+��W�;��O|j�R}�4��[.8�bO(rӺj����S[N��t��O�M*rs�ʖ'"��Y��[���%WSD(��uocqg�L��THP��ia$3���ֱ݃BI�n��H!^�㮓$HI����iP�$��sBx��{1����{ϛ������}��gR���k���7����ti����N�X�� v����3��@��������E$��e����Ԇ#zY��=
�8܏d���[
�?�D��mY&��dD��4��ob�ί����rHx��aC~ӯ|Sw�eq1�~Yg>��uMy��׾�,��lI/�6f�G���I�Gdw�����z^����w��mM�r��T74���u>�}�o��	���X����Z�9�SǪq���V  � �cj���;dqݕ�g����q�hA�K�`�\����i �Q�V�;�������04d�X]/��I9�x�ZK�w�	����&��@�k��$�>8���P���;�{��b���8����0��+B�.�`�<_�I��}�{�9O���7Y³�/�8A��u��)�p����2[�|ۛ�A�Vɒ)z�SL�<�;�� N�G(1rp`��8����Z_�jw��*Y4i'���Y3j:��/��$�-�#*�� ��M#��޿0��7��[����)��W)O�h2�|n~0�|��Q������R�^r1�~79�,g��O	�ykVL'��c�ύ%#A�	z0vF�Iix�392�κ��W�;M�d9���4fHX�x����Ɲ���L��9�q���F���v$CSO�+�����;3K�6X^O�v�ӷ���E�b��א��8�աc�OOlVϭI�,�	'C�5��߇J��2(���e�͞��:_�r��l؇�I�Qg��,�3 ]J=���
��UƏ<��xټ�f�IJ����R�d7��9ږ���h{��δ$�SdK��<�*�"�S"�A\�e򛂖/�3^ h��+:�6��#u�㾱�y��m#��V��Ұs��?mlsv �t>sQ�՚F�ޗX�/7�;�P�<>�w�	��e�&��H%{/������(��B�__X:��ಌ��0��xȕ$�cI����bJ�z����Ç3�k ?}�[�@΢P���fe�?�*�@���R�Gw�.e��RE@�(��f��9�S̻W1���}y�Y
Q�xp�:���:ڌ�_�m�'��_^�i����Ѫ!��n�[6��?�
��H�j4��5�?�� |����7,}�ʡ�ћ���E�or?<2�����SQ�=$	���.�cT{�{�~�X@Z��Q�)���E�-dO���X%��x�W��<���n0p�$7�c(?��c�����}`�M�_^���Y{ �ɲ�V����֔��V�c�[����%�]cM���7��U\^&rZ�><��X�$��V6~�k�m�{���I:L@f������V���	JC[[x��B9��7-�q)+����g��;�PƊ� l{3��^�yo���m�!��8�Ɵ|v<�4 ĭ(���*Wߑ�dnT��Lf���5��++.�����oR��:�þʢn���0l��[���͏�/V���w���6gx�m�	&��y�[����k���>�g��a�������D�1Ϊ�0�?�j��n�Qf�w3�ʮ��!2%Xէ$��2 N�$X,�����[G܍�W粆��#��o��J�ܶ��Fv�R6UE%�3��<����0e����m�y�U�Y���P���@�{�!{�z:N�@F�9g�H=����;�]���(<�����N�Ge4bQ�I�����5�/�H�ۘ��A��Q�h��@+�T��v��wE��f�5��-S(�`��r0����8�$J�%��!�*���S\M�5:�{pww�w��\�݂$�;�݃Kp�!��������?�V�S�JR3�{�����9ӃG=|� ��q� :�NǛ����Fc0�f��>$9#J_䪼� ����9�jғo�M[H[�L���>ETs��Q�~> l,-���/d` ����"�oкՂ�,4���#�>9~� �Ȩ��mк�6�ҶF{[��K[�/��G���ɭ��&+�N�E��yL#F��r���R݉'4��&�j���}iz���sił���3�G�. vѯ�?!�����Bf���Z��{W�����z���:Y�t���p7A����z�1�8�&ǩ��t{c
�U��g
���.16�0��Ve�����4wH ��#O~��u���F�k��ل?����p�g���1�՜�_$!_�?`���6���[-x��d�z�ST(��%^U�9�&�Lw��Q��1�����&�:*=����������WO��exPv�l��ޗ�CT���xs�op7򴞝�U����M�x�~�z1�����JXFދb�'����Z$�t�=�`]�}RwG/�;��>o-���)ԠyY{�]�LY���ވ�R=\�0ZKV�{mkί�o'�c$6"|YJG�V��[��Nb�L��B�sV�����˿5[7�E_�G�`B؟io�(���~n�;Ǥ� Y�'���~�Wѩ��֒u�R�|��i띔�D(h��C3��/O"D�A��ƀ�5�Q�PzS)�`��	�<��\!�K�p���^�m� �Sv��ń�^g�N:#F
�jy��;W�%�q���X8�&#G�@x�F֖ݟ�O�Xx�V~Ub$�h�z-I"�$?{}�x4qLˎY�IC���̪A�h��<���ѝ���	��q������i��2`B�h�1&ˎ�笖?u�*�E��!*�Bd���J�W%��ʬ���=����lR_��ڴd)��~{��!��u} ����S�ma7Tj�́<�F��d��l���IOJ̄����;�6�:��Q��,��S��Uo��<�6�~�	L�{J������UI�g˷�qId��_п�¼'��`)�����!�u�K5V<i�����m�!n�������J�ۛ:�(�.=_�G*8��E����rj<Z�5���6xr��iNѠt�SҪ�����&��~֪���{�F�P���Ni�Ռ�^�G���Y�ӪD��r�z!� ����D$8I��Q��mKY�N�-�B��ā�V��\$�<9�̫_��C-T�5�'�BYao�޻�͸}^��x�{Pw}�*}�t�T���N�L���Z�����E���*m�7�����ᤵN�)w&����{�}��;fU����6�%\��9\6�Dt���b����j-�.:�2�V��P�F������<g����)�A�!\����ϔN�\���`ժ뢥���4:�9��G����/JbD�cbH�&P��W���D	Ŗ���JJ�\�F�F�I��-Z����J��I�k f;�Mo��>!y�`���TLf�>'�94h�lP������E;��gT�"yf���J�z�/����)�N�du�7�����;�YFX~��R�҈���4&��nq��T!3smv&zf�����:ܾ>�lJ��JEc���<s\���<'�����H���xc�
s
�Tm��$X�0D��;���&�Vs��?��$%�lV:a&����>sb=��=z�D#�Yj:�d+�S�o�~���3��;�,C�"b
�]|x��e蒗���%�� EƂY���	>Y���a�e�Ņd�6����7�g�^#_�����t��m��[M�Q=���A��	zOe���4�V_T���3{�i��4wC��Z�"э@`_
�Y0�tur��?Y�<Y�֖g�L����zy9I$��/��F�9�����d����%lxNo�=����W�T�M�ǎ���h�1��@ҨR_��f	�61����y���=-�?�&��rV�h��*�K�:�,�^?|M2�mM�� �V9v��ѫ�*`Dr�������yz��Y.�Y�W��x�&��9�w�0K�ռ2\w�nH4q�Y��
$'����(Z�V�"QG��2Z�5Ԕ��O4Hw�x^��LZ��I\JRz$VR��:�����&���������]�����qfT�(��$H�Uڤ!rн7�A�X�Q�۷+�����Rj�đ��>��H~Z��e�`��<`X 9%�~��? ɾg*���S��H�*w]J�ND���I����'�m�)��A9ip��JL�h�Ĉ�����%>�y@@:�4/���r3@	���\+D�-�D[y��溉;���Ut�9Żp0ɵ��R�A�S��ʠY�����]k�ߍ���w��.�,Wä��g�ǚ{~=����Tۃ���h՜�>L1��.��B�l`$��5D~L��F �w��)]z�3/Q�����\��*
$2�n�*q5(�4S���|�2�Q���SX<���
@g�OU_������9�����G1o�wp�u�&iC}�ar�b���L�wT�1�Ñ���t��ް��c%O�~)���x�>����s�F%�*�uĹ�	��(���=��}I�MFy��Jͬ�A*�,W?�����-]��$��'�$�l���k �e]J�1�rVl��w ���a&f���ǃQ��d+Wĉ[�V�ɽ��:j_�������}���x�"���ϒa��F�48�Л�"Lv�6ō(!��������}-<��,�×������3&l
�j����OY��0��o枾�iYSY���hm����uѦ��G|�1�+�1�A��y���Gg.���,��N��=c�S4PP�1�3I�����ͥ蒡�]�r;� ��z̲�4�uF{�~Z*܀b�np�"P<'���'��R����e��	P��O8������W˃N뜺����ä���Q���_��m�7�#�lf|�&v	I�%����Z����)��N�!��sn�D�rS����Z,��"��:?�`j bh�k}RL��>��b�&������mj��sy���9�z,�"+�7���12,�K��-@�ϤM��Ҭ�
�bx�%�W� ��P.��4��=�؏��@I���Ь�x(-��眄[6��F2+����Q8����YaAlC�\�L\"�=/�w9���Ttdz�ɉN� ���Ҥ��4.{1J���'w=_���5E���Nw<!��f����G�k�j!���2ǒ
�Ӹ4Z�_(�]N��
 G��+QN���y�X�O�!�\�2V#5N&_�іo�0 |�NEl��Y��4�$��!�*��
�b	3�����P��G�v��_�!��͵tA���/�/�y���k^��:
%�T�J��.�h�z��Xڄ�#\�U�7�i�ʵ����J ��m@���U�e	���n�I��;���z�}*��s$�º�La)��� ���|ǩ�#@z:x��}�ϸcZ��LB�Z��iZ��2D̉�^L
hOd���b$�
����HU#����d�tW�.�4���ezسY���I:����S���ضke�(��a/���1oj�]XV��g-K�_ِ|���D*�Ts� G��f���Ӭ����_��'�֫#O�za���.�h�|)�0Qr�g�K��Yx�E�ӖVd;Y�s`�aRhA����AZ�c;ЮV�#eD�o�J�+�|zʨ��Ө����*�3*N����L��=���Բf�aY��نɋ����Z趣,�ɥ��OMȁZd��m���c����tBׯ�F��p����Y�q���z�(wV�O^���+���Xޣ0˖=��z��g���6>J֮`9��E�qU  M�E
?�I�2��yO�T���m���(� ��r`gk)�Y�H�j���ȳlB��^`q�y_��ih�-WCa�A�	�z�qav�*���qj��v�DS��Ng�h$�� F_��^��6���r1tvtY�	P�3�	�z8�{�
�ś�c�q���ì�(�\�=T\A��t��O�L��?�d���?R[�3@Ub��)��R<�S0�(����%�g���Y���IC*i�lד�Z�V�Q����5I͌U>}��9/4�#�l�c]jl�{��%34�P^�E��u�����cY�V���a%�ƃ?��8��'�RF�;Яi�^/º�m�zg]�Ty.h�sb#�J�Ԝ�w��d5�>��uka�O�I\�崂���ia�4]kζ�'t�%��A�r=���(mX�	�ș�o�0��7&��(սb[�� 8���0Å�o���|2��8w��=��)kD��I�ŋ�d�����I#+��ݽ��e�����k	�͏�@ar6U�a��x�ìv����iC�� _.;�9(n��Y�ʧp]��Οk�����6kPh�"���V���:/Z��i�km�G!P3XX�C+�{�Ї`ghh~�d9�
a��%�q���?NR%W���1;8���%��A�����W��������x�e�@�C(��k�a�+��+����d|F�f�LO����Pg7}���-��èF/�FF�_Ү����nis�9QY�f��M|��� ���Za��G{����4����y&C�kmM��4�gF�iZ̮�k�V�Ƌ��7��X�4�������	J#¿C�������1����:�Y�<��P�7��O9���׺I�9(C�0���vF��
��$�}�8y.�����3?3��٠,�ph�Y=-IrԳ�5Z2\�#���6����>�����{��#Ɏ_ln�@�R����h3�?���_��[l}�X$9�������o��=מJ(˔7^2�>m��/��ԿV"I|gv~/@z�? ��ME�b���h�"t��P<���`y����ꃊ�w���e��R.���ŷdmkd��  �&���.�	'
2�b���L�{ꌧ�Y���L�7�(�ZpX��%����p�������f!����a�����O�/�����8�h�ߘ�Ja�|�ʗʷ��s�t�f�܅j^X�)y������NHr�<h2�!�w�+b(LDG�%�{Y͔[��~�p�\�2_�:%�E��r�S��lQ7*zC�B�����&�^��G����q����0�Fz��7�F)w��0l�GY`���z�R�@_�M�0�S;�����5Kȣ:�òtK��;�h<0�Y�S,�U ��(�x��P�&W����>r�mVE�ᨖe��f�;_���Y�.1�����R1A���l���G���|�as���[���h|�(�ը��܇�\׎��s�sB�9�]�\bS�l0pWf{�}��"� dF{�G�]\���~�N��#c�����Q���e��*��z��w���D5uE��f]=�W���6�9Y{�jo@C�8����������)з�:jg΀U�;��٫�î�
���ӈ=F����$.� �Eq��[�������ˬ=��0<��O�&��-�׳��7��w�z<XI�������:�@�Cݠ\KO����:���b�g����QO��c�8=@1�Š�.�H�[["ӧ\�����Xq]\&��w��Zw��7U&�����^0�xK0�'<�c�g��0*T��,�9��ݛ�P�4Σ��"玺���(�"�'�f/0Ѽ��M�B��p4��<���iR�����
�a���ﰝ$%�Q��.4���*�3�H��/?�ԄI���5�y
<��!�֕�;F�4���D�,A��FK'B'��S-�������>�ǁ��韗�T+����t)=V�S(G]	ͮ��+���4p��֐nB�X������n}ģ�5�J�Y���$E�������}�4����D�t�Mo̪5.��o�	l+/m4�)�����*�o����Y��P�'��$dJ�M��	�e�jN�x9ܝ=�|�QB��zQa�˂LL������c1��O�����`H�-|Ș:���p5�������}(���V��<o���D��@�n�|l�ykRв�bz��[
��'ʹi�=I^I��HV��J�ne�9y'r4�ލT�D�D�h���a<p�[Zz��Me��Q����]��{�O:��NφEX��ʺ��Yǂ����Ig���N�T�'��?V��������=��0A�;I��!U�{���/�^�d���2��r��	[���<���G�U@�i�A_;s�EyrVh��k^K��x`�?����:JF�:P~m8��`0��u��d�/8�a�ۨS�&@㫞���F����7��r��d�^�bҴ�!�,�3V�	!�w�
U�B!SL9��p��`��a�����i|��]���v�ߛ�P7�%�B���d�ϐ���s�A�8�c=�Y��ň�]:ģ3/�&o��0,�|�5�_�x��1h���<��+j�؅͠�,o�-��B���cC2N�B,���%�)ȅ��p�����FOv�s�:G.���I\�phYH�f2v�0��D�W�l�V��Mq�`؏ߍ$�n�/�W��>i���	�ϫ���R�?z��؜�[/�gx��ġ�v*�:ѐ�Y�k!t��B����u���l˖�h�s�5b�F�J��*ҟ�i��g|��c��ײ��Z��h~�<�<�;�����1�[�m4T83�""�h�i�'�#�{GW;�����G:�+mZ V��T�����׻]3	��ĺTZ�N�2�d"F&T�S���1��� ���r���=c��xQ��d|��i�z��hGt��Hd���V�M���l�հ���������K��C�.c�C�T��0��Yy�6R.��$����&��Bs�D�Z_��"��ڐ��)3;廉o,PS���T =�	 'L�.�k�Ǧ��:��\t�v�V�Hg/G.��ځ�&/�h��� ����J����`xQ9�F++<�xc�{��懎{�ጓ�!���=��u�ߋ�����,�Gl���CM���L�m�5G���q�m����`�Ţ6�He1A�I�6U��@p �j��/��MV���G�c����N�1�h����)%��9�no�coR]���@�xR���\��j��}޳��rW#e8����z�W=o�6�Y'�����[`N��P�x~xI�����Y]-G:O�~u�_Lm�o�Xќ�b��������	���
����P2���������\3�<#S�Jj��d�EyC{ĊwW��'K���e������(��?���V ��/]]u��v��ygy]�'���O*����q;#Qv���'���]����d�v(���g f�>��"�[�ל��!��d�l1��d[e�&�OQ�
�g[Ggm��T�(����̹~��;��cf�GO���-8��a���w��(6����_,����R�<�P�a�<��d��Qn�=�@&3�G5+}�2�B�n��Fط� @凮\\��U��!1b	8CUd��Oa�|.<<8A��o���q�(��\�:\^��>$���|]��N��qSqq��#s}�PP�x.+�b|�~3G����KA��+Z�G/w6��B�CR���&��d�}O$�Ǧ�i(�z�@��F�V�b)�'�i�C��*�������F�j"�:�!(!f@a\�1��O�) t54R�B��B��,{nB�u���3�/�t�2�gǐچ����z�@�:��=<|�k��{�SL*C��uz�l<��d��ly���y.�Oٽ�&�GL�gm��@f��p�Z�b��&a�؉K!��JʕB�\!8|MTG��-w��w�(�`rm҂�_wk���A1hb_�WP�����'��3��O�GMt����>�@����;��*f~d�g�j���P�-�Xҩ}s�M-&��@����$̠��4L�Z>����G���[������H#2f���f/܃�r)��THuH����H��<�:pzT��[���XVRd�NIm�6�Y<E5+����s�U��f���Ay';���l��H)
&����\p%��L6o��F֩����m~sd�Ќ��F��fy�ͩ�p�����͝Hڻ�޻���m��o��p��p�t� #_�?�U����������<��PU%4�>�����R��^��Q��;���[���X>�3¿R�oV��z��F/,lV6�?�Q�S��J>[_���#�N�(����nJIn��K8��	c��b���ħƉ������/$a��/M#zOҨry+�w�a�4pf��~�7��9!)��8n����S����l�8Ӷ�n6� �\:!-mA��v�T(8��4i9�dBB��QGb�b���e�.�w��kq2�}#B�b��׊�Ȓj����q�&�GB�o�e$�Y�������S[P<�Sš��9�J�����u9�n�⦾�(����<�
e�����gb-2��l'�P�5'�p|�Nڷ���]�c+���wm��
�M�1�u�;�v#�U�ț��%���.\JԦy�݇����5�%#dy�e��F����a/���>�cnǂ���>�q*��
B�,	}3���ϱ�1M9GSegɡPH�[�U�\ew:*}�Ж��� jM~��+�ά���
���P��p�Y��&�"E@>���f���1(�Y>��6Ծ���{�>���)�e�ba]��@��D�����%J�DJ�]Ҩ�����>��4�h�M 
�dL��b�.�����Z wH����;��.٫���5�|J��J�;z�c�d�l6�7g_e��0R*�3B�+(�*Q�"��Ai"s�Z�)�g��C��S��Ak�R�x��x��l�!�U"=���w�5{�����֎%��5�V�(8� ���;�=8�6l#I�f�	�s���B�|>�2. �͍�C/3i��P֒�˹�QiX������zO�cq-�++滘�~��D�)�T�`�J�������%�C� ���,�P�9�l[I�!ې���7p���)�Ȍ�&����`8���Z����n~�� [�_�
�Em��Q��<U)��Q�R��Qr"QZ��h"�Gj��.��
��0=T���h�yB�KTow���~<�QŻ���*�ʋw,�����$�;$�]^J�P�|�s�πds�X��1��>e�(����n��h0���B&�F���煄�z�'zv�k(?H;����w܆+4B��2��	�}W9��6����5�6�8�/-�9%T(%4��B��e�����N�C�^����s�	��$�r�7���R�^CL���.t�8�-�-�\S1&U��ʑ���%��3��M�`���Y]Ht�& RtS?���4�ݽ~��ZO��\c� }�eC+��\~1GŻ� ]�a\�+:9k�v��\(�`���4��֒�d�,bZ�6t�bdK��w�	I�tFW�$=���=15�0X��]/�;�eQB���V���~.:%��k�[F;�Ѥ8�5]���߸�.lt�����t�q"%�CD�CN�>�n�t��晕�`v����������e��ZFq�qpao�j@���?P�%@�S&��Âz3��d���3�ϖ�9�0Z��+\hX�(P����[�h�!��E����6�e�;n�����r��e�� 1�Op%CO�2yT���V{J8�����v�oѮ"�Rb�V�s��_�u��R�"ǋp�C�NST��Ȃ>�n�U顋,9F�%�˨[J��_�_����w� ��ø�~��!��b�����Bh�Z��|<A�@��s���b�~8,_3=Sf,���"�N�f�S����9f�-i�w��8FS.�_�xx��ۆ�.4�	f��6Au���n\%�=��;,TW��EG�L`Iɜ#)�ՂY�����.bȈ�����X����3���`s��ȩ�H�%�����ٳ5I�j_ś�]XkQ�0(+��9FaCN�T�����rm2�
ra9$[�ѺϏ�s���q�z0~N���X��&��a���SʿxBrܴo_N9 �n�	�d��J��o4,�,�17c� ��a ��� �w�D��M�;Ƣ�b��Śk鱯/s�8$_v�`���W?� �%"�/���`8�~+~
���ڤ�Ʋ�/�'"��y3�<����r8�'.�^���k��b���ˢ�~j`��"�K����F-���Y��9DB|>m�d��|#,��sG���<�?+0���)���@V�+�.��
xKV�r����ixmt,����B)���=��/]�itM>/�ɐG�$�7��7(^^}[��{�id�.wPU+�dY���]�i$��/�2r��>A�ӐA(���*��m��tòBN=����	���_�?�E���tDS��.�u=�Z@�/�ѥ�?�g!]l�-/�� ����atx�������?RQ�ߦ�<����A��;�C6�tB@���H�[��~�,D�X�4���_82���s��r-T���*T$_OI�{u^n1_$qw+y��0Ch�O��1��Y�օH�|i(��mA6�]���mif�_���N���f�RY���f���~0{.��;0��c��{c-��
��\k4����2�j�(� ��9>p�p��G4��D[6���0��K#��D�yu���?u@��J�i��V�d�n:v,�;ϫ�������@iL \���(}���Ŕ��;φ��I�s�m⠙jfw->.>����>ϫ���٢��}�>>|�	�- �P��k�4������E�� BIӝ��pZƋ=;���2=$�{��� �ẉi��M�.��Y)9��EZf#�%P�����$Q=�bc͞���\E��G3����e�^��\�c�sF� �ܲW���T@�sK~�~^�e� 4����}���n��݈o81`+� V�_�|Iu2 �ZΈ�ͭ"yI������V"��p'��	�0{��s���].�3�j⋞��y�u~��d�?��&1�		��V���+�j��m+}a��h@P��EV�7Oi��k����村S�-L�5#:��� G�E�2�FY�fl"&���W��V$zG�����u>X�gß+���dd��-q ������ͣ��p���Ķ圜 G���'��c�R�Ԇ\�"܌z�VtLk5�iV���{چTr{���Jg��B�J��o�'�ͺ*�����g���r(��`d�kvV���B
���<��,��ZYRO ��H�ʰ�����|R��}�-[G*b�{J�p"��:tw�
���Au`�L�wз恩z:Ծ�
���'�g�X6f�<�*�q���h>=�]�;��c�弳ʩ����4������`�����W�V���m L�V�sB���p�;ܦw��5�w�mWx٘e�Mߝ��4�H+�~�l�I0���?fC�ܴ�F�S]'��#��ί�gy��D��ߨ�q�g�����Ε���$N	}� �f��X���2p駫�_��Pj���ըO�cI]�����cjm�_���(n���C��'���AǱ��=x�����S�1��k�n��u�5
�k��d��i��ýNJ�,{?�����z�8ıT� �x�!�@���X*��	�lgƏ�9�n���@2X@T&�p+2b�Z��E��E��g�+8�}#�Ȩ@g�l�{̸�<A�����ʹuf
s�t���C�-S��]�W���!`�;���@\�#2	v%J-Q>��0 i7Z�j�R����\҇ќՒ�hO�>|���<��M��c�4B��Xj��	Yu��6���%��J��?���08_`QD���9j+�a��d���
ȀN[.d��OTvљ-`��o��p2X�u8	�^N�ve@�q�i�ri�%�1�H} �hցb/�6u���Rse��p��ć��v�I�E�@1�!G:	(�7zt?�i ��c�=�+/j$	�]����ʖ��gϑ)��n�796v��$b->I4����nGi�il�4N���WU�P�)]H)GW�;���'=K�HӤ9Dc˟յ��C��>����Q뙄IK��)pꑊ3m�����U#ʑ��!҆�(=V<���W,{���1u�#�+W��#ԭ#��T���@�S�s�*`���V�5�keB��{Zԕ�rK�kH�[�*��y{e{e],���p�v�)��v�ϑz�p�����a�a�Ȧ�-�T��RL�~�����C�0��P��`���<�9nd_����-��i|	@��	������{��04��~%(���W�@�m�^5���cq�� α��HF��9�sdtN��^2]q��gN �)_K����.RX�D�%C{����S��4�h+	o`���D �c.X�>lVFM����2�N+~���ч��|J�@���fE�������+����_���Q������s���^��p�������~���{%#���^篒�/u�����OL�T�9�{a��׾}XHs�L�j<[� ��-�"Ɂ$�%�GM�Ź�mp�l%�k\�г+$�.=���sF�o�q�i�����Y��[��
�����TM�����I���6�3m"���"�c&$'	�^d��D��W�R�^R�Q��$�
$�����|>k<����9��T��4Y�E�%����֠�4���.�l�Q چ�	P-���#�����\Zq��ow`8�l� X�$���|�ب@ι��^ތ�Y�\I^=� /)��C���c� �|~����p���+�dԺ��7w�<��x����8��k�␍/�Q9��i�zf�h�U��/�N��� �Ow�o�S�-����?V���:6��S���s9�`"�
��Ȧ�?��V@�\q������rG���l ��b��u�����b����!S{V��X(ן�ѾL����b!j�9�A������0��8r�{�j�Ѥ�NB�N:�$�u�%syv��
>��� �)����JF�ϖ)�!.�:>�8�f���� �}��TwA$(���?����~�]��q�h}�$���q~�T�>A�~ڐV��L����p�UR~�����w�c9�ȭ�'T �cH<t��2����q�d�@Y��2�b�n�ÆV�ъ9d�n���gCOha�AԾ~���t��2{�n¶�F��_%�*�J�o�O��.�I�gOG�	��i!lOc����x#b��A��_TF��E3�-kz�/��}���?�yTä�~_��72F5L�����z�=�J��XD���2�N�<ړ�;�F�0@ˤ��� �&g���!X�n��OT��W�6da��η�ߑ�h��a���ŭ��q�\�ӫy�U	bw�k�Nu�a�75��ٔ�DZ��x�D -}��ҭ�d,����d�Pa���?]]� ����[C>r1��1�
����~0sh�v_������BTۑ��$��|"İ�I�N<�Y�/�o�7���l_���!�#���E\��)��������f
�D��j���!����>�<q�A���uSX�ݦ��#��c��}�xCx)C��6����ዉ�����Ą��Ro� I��t�1w���[F*����������I�`T�
�G�E�t2QXr��,�(���^�L��*��,�z��N�B���k�˒���=����a�R�7u���+���H�N]�oI��Q.��N��
��Qs|��ۛ���J��l�s��g���\�@�'Mu3�h�Ê#�77IYx��&��
�0E
���ZT;��w��?�wS���XXz�:�H�UYNkm(Y+�
��.�3"a�TOd���'�~�۝�������J�u[�1����%/��1n,�v�V�;"n�z��}B��E,)-���u��rҎK2Kd7��R��A���=�x�N��T��8�Z���Ͷ��u[L���-N-*�J�XS0�Mo�C�*�$�+|櫖Y�g�S����]���Ni�r��n������%Z��wӒ��W�/�����#pWb��|�\��������w��Я������B��f'(|u�"S DN�3tz�X�`�����w��y{�o౦�N���Pw��Q�.���*��b��u��Ch}B��$��Bx����l��0c��@9��y;n.%	�OE�>��\���ˑ��S8�AZ:Tuv��p����5��1w�
�����Ƌl�(H�b_7Ҕn������&�;�u�H�V$�E���3�ڇge�rҁ.X��b�֢`k�]u*�@��N8WZ<��Җ�͔�Þ���C�1�I�I�u�OC'���ڼ;}�&�O����ԧ6����W2���/Ɲ�KMW6՚����NCv��@�I���ox:J0�|�`ȹ,fP �E��!a~_W_z���s��,r���w!�A{0�?��G�Г�o��g��Ͽn{���Ճ.LYG㸮�/��ˀ4��rř��-)�F���_�(z-��Z,8�uƮ|�eE5�XG�ɏ�M�K��-��|N�������Ssn��Λ�����e<��0@]����{��A	|�D�J�(�R��$Y���A�Q�N[�"m���󦁓�n� �l5O��VƯ仚��C�:ּ�oM�z�d���͵�Vr���jb�輩�Ob��F��&���%��,���Zi�yC&=b-
��NҝD#f��u���ڇ���k�t�c��N�}��8�Z"��ƚ�5�y�l�C�N���E��|����ޗ����T�����?s^�=;b-����0&�b���l��W�qP���q�&fuL���0egA�)�q�;���Z?���%s]A+/������rq���-U�C�4��&��#9��8����e�(��ۚ�=9n��$q.\�$�����Y�蔃O0��z�u��ތ�:/G��A�t:��������@;��I	�a������ed��YIۥ��{z�ss���ihİ�4E@O�w�AO�\U$"����K��I��M��T������[pF�g%<��>AX'��߉��X��fQ�s�}_MFґt�/-���
��\�e�~^9�����D��Q�����^Av���c�x�g�ΛU�-g?�s�4�3i��p{��r9�cg3ҧ�%�!e� ��Ibs���@�t�����#yL�İ46WR`f����Q~!�>U�@'����J��֒�[��M_��K�����5	��ᤛI�)�Ck�p�B��Q.$����ߚ�fe�&(U�o�������S�4��k���d��;�W���^~�7wt��6�l�K��qYWWX��u���Q�y���;S7x�{��������Y���<�w%熪f��&ߘ��P"���� RL���Q_U�T{F�Q��	�IE��շ'�n�#R�Q��{B4q;x��
��N���Ţ�]�Zh1y40"ֿ6&�]�D�U%.�X{��=m��*�k���Xp�#%f"��d۾�܆d}D Q�;kCGN��H',1������S|�ъb���A�A��*�C��o��\+�d���b�7)O�qJ�Y�|$���O�c�6��T��1C�{����1@x�������M��⋘�!��{5ڣ@��{_m[m��UK�bOTX9D^�@L9�ae9
��K?�O�ʟ�2$���D��	P��ORi+u��m2o�Y4�3��ߌ��ܯ��Q�̼˩m�t�;\脐����w�q��D�����?��8F�WX��{9ac�5[�	%"X#��^Z��BQ�
�7��{������4�]s���7<��+߾%	h�O�ZS[�ݠ�{�c�y�7��ew%6?�3�#�!RR��!�A�ӆ�J�&�>E1�iy~�����g������������5	�z�Z�#��n�`��������UW���Ӧ�|Of;A����{�`��4h87� ����4��"�k�k~���f�� �_���/Ә�E�y��ws��t\�O�Df�W�pmYJ*���T�ާ���83".l��<��v1*co9w��b���^{�9z��[�-��GQr�]��!�bWo��Tɽ�3S��EjhfM�2^$k�Ҽy��|Ж���\�.�ϊ�nN^����o��Κ��a���a"�C�����Ԩ�UΆ�4�5Hl�Z�O�$�-�٧�90�Ȁ*���WXU�E��&�~������_�+d�_i����~�>�toA��Va��#���h�!��{W+Tv`A�q��ih�V��M�A4�PH���O��fb�!Ϟ��).�Po�`����'����QL�"��w��Dc��ֆ�[&�:���V��ڹ�<�/J<ٿ'7�c�'��¾&����=)���`^p4s���<�JF�#l�IY���ÒY��0�N��ݵ*k�(��f&�m��"�m&>TM��\�v`�X�U�������aE�Mȧ��K4f���=Mp�C��.�1�C�����@V����V��_b��g�P> q\Х��`W����a�]��iC1A�wp>�^g�bo�A���"�gV4'TY��7�j;a�ȑ���#�9}��Tm���=A�ϼ,F86ٚ1Ȍ�,��C��=K�2C>�c��b�0Fi����j�3_�!�4C�=U\�Ch{���'{�+E^�e�MO���hh8�^ؤ��X�<r���∅&2b�R��:/C�4����<���c���B9OZ}OI	�)�����4ϋҭ��~�L֮�s?������%�	;6��sg�?X!���s(Z�f���ܢC^�������$ZE0z��3/lF͂�'ē�-�>w)��إ�����`�?���>e6*J��|~j<�9�(�`��3�y�Tż�5	���+�
�Ӝ_˜&�O���<�
<	@�p�����i\������������i���Bb�l�[�渭xk�E?ִX�=Y���ώr��������Z�Hɷ��s���>��?\}u@U�����Cꒂ���E:%�K��A@BJ�J#���tJ#)ҩt���>���?{fwg>S{f��"�]U�d���{J��ّ��ٵ���ϕ���^�a�{č(�H��u,��c�O>�i�Y�����;g���|���5��8y�@�.^r��.���5�y�9���冟Yi*c'֤���b��^,�C
D�J����k���\���:���ƭ:]μ�73oYeR8CkN��s6d�1Wfy��_�y�:d��Sq�}>;(O��eӶ���FQ6+�z�C��Do���r�l�\�~[EJШ��#]�P���<v��-���},QԒ�������?*�W}}N�7� �L��/�k���Ifa���r=�ߐ74]�+��%'���O:SF�v���"��� kƩ!
�<�����.�S�Y��z��&�'+s���/�~b�����W&�N�y���"��&1�t[\� ��{��g	'٦��Û5��ד-�@*�1��px�h5�Yޤ�ў���z+���$s*baR��|�B��<�Y&7.��E��y��WK��_�_��	+��������*���̹"U��m��)%�.y�7�.T��� [��|��@������J��+0�c�>�t�J2&rȳ�K���`mN�O��ҋ�<w��v��\_���J�
Pv����N�t8CZU��J�a����-�L������r:��#�, �˖ok��d t�����VdfSғ�*<f>���?c�"�rC��������{�[�%6��Zh��X��°�2��:�!�喯Z�(��+I�}> S�)k�.2s��L�c�1��ę	R�7���__J&o`&���o��+k�K��r��t&<|Z�����$v��GD���k��qf
:����^8}�U��m��jS���^�f�[@�� , zϙ6��Y�h������ֵ� ��H˖{������-ky)��,|���e^�|�Z_�%��ن}��o�	�XT����{�¨i�b�m�����q���\s?�ٱ�~K��*��1����q��x�Gd"FY�`����	�`��BT�]=F��7�'3����b�p!��b}G��];��m�B޻|/_�˰g�uq�!&%��wC�H���4�oVx�8���tnؐ�yx��y�5,���Y��M�z��Y���0S��T�b�������F?>A�u%���h^���nm~�v����R3���d���{�jp������� �,cQĪ��n��O1�.�E�#����~�6�}wfF����.1�;g&���y<���?����fSج����/V1�U:���.��G:X>������>�^oI���Mx{"�˾���Љ���=u�a�n}�(tALI��!|�w�s��<h�t|�;l]x���ru��<�f$�����ކ넋ll���z�J\�=�T�.����*�J��K�%U���fz��d��~�X�y��u-��g˅�kz�d}�ϭ6���w�s��T>]Rݬ�Ni_yH{������ɿOp=��G�Q�t��ryG[d\�n��>Kyu��,��)r��wl�n\p���J�fi�ތ��XՖ�-r�Đ��`L ���! AeߤБP��l��7��Lfi|�)AX��-Ҷ�g�L�8�ӣ|,�?/C3����Fp�O#P��H�ʢ��}eB���^ � L�L�� ��l��N	��5Nr���=��m"��s�Y7 >�\d�?ʶl�<ߩ�f��֩W3�	���]7�N֦u��&��@�(�Q���;�.�vV3~+���Z�i+� ��5��O��ܘf��bKXr:HI��BY��t����4z���T����˦'i�8�|�
�37aX����羬�R�7�a�}/H'��s�����О�J*�|����該��=�*��/l���I|O��ZQ|�L�ʅ�+��-�~Sv�Q�&g��H��)�}�sr?k�A<"�[��RBZk���>�N[�/	6">�X��Y�+$Z*�WJ*�T(��C�Ƽ���I������՞VgVm�/_��;����7��լ��g�����}�	���:�V��p�%䢟��K���_��'ۛn�bMJ���e]^b*��6�!��'	5\p��3|,-��dZA�S�GWp}�~���U�G�O%�2�����dd�bS�s\!bqqKq�:���m|��T����������-�,�_!�8v�\d��w�d�p��ҀO���D>w��5��
*6�c��օ7�>b#�����.����]n��[�V�m���!u_�`�.�%��#v�u����{��%�����54D!��DF�ؼ������ٝ��Q[�g���RRZs1���f�"��?=�F��VOP~�K8B�\�򎂪FR�ng�^!hSt.^&�p���~�����������Z�t��U7�*v���̾�f#�-����y�u6 �0]�n���K1q�����S���*����N��@>����HK~�������3��mpK���җa?K7��8��_����=�m�k_�A�2������X8��.�)|Wh��*r[�s@N.��V������.�hx��7=��k��G�1�D<V�y,?�f�b7���e���΄1�kv��ջ~�$�興:�P���R!��<�&��A�9Ӻ{�uZ�Vo}�"�;G	�NE��d�Xpy�5��o:�R�	x�wib*�Vp�d���na�V�(�.��j�O�L=d�qpR{��_�E�����*��˨< \��
Eq� �RBW�6��v�2r49E'n��}^/3(��CW���N8���T���#��l�0捍��	�ʬU�6�6��T���zE��fI��kA�sB06�rcB<��I��[���1�;�E���ḍcX�¶	4�8�~��RWy�4�}fJ�ź9��ơ��ݨZC>�h6�Yޟ��Z\?V�}��SǞ����\��~��" ������|��k�:���Ͼ�����w�=k�J�}^�4�NΕ��ϵ��g4�rwRJ�k݈[F۷:�<�WLR!-+X���Ǽzb��	�R}�u�/�9v�{�M	!J��ɦ�{�M�Y&Ɣ�b;A.a2�f�YTe�3сP�_Q�����h�����������=��e�ğp�B���6����L������Ul�3(fB �r�����I�jB�`i��f��C_k�d�^6��ui�=�h�ρ��Ѐ^�-�=��D0wNC!8�`R�bC�I*��� F�Iit�W0O��T���sW��+��'���m"h2ڼ�^o��l����D]�ÈMMpc�1�WDLe��7잌�8�tmF4xZ޴x��i��'��� ��Y-�!�\�^��!��D}�㙹����t�ݧ,e�5��A�=���xl� �R�{�$o��{V�q�,zt*o���7���ڔ�����ªz=�'6E>pDQ�1dS�����s�]N�׺��z!����L`��
�f����4-�)��sO��X5���X�t�VppЈ��7>��U���V��9I������sz�B���B�DS�r`+vm��"OmE����D�2#{hZ���k����TK�	������+Q����H�����x��􏮺/��j;�?�ʘ�b����U7�0W����&J������ZP'����=(������4>>-ٲ..�̘�0�M�&�%�c5F	K������c�̟�tӘ�E{Q³��	_�BS�y<锦��#��5���GgZ�|\��:��Ѻ9%� ���B���h�1���v���*�I��?�i��7y�N.�A����/؞zv<�)�<3a�f!n��syM6�͞�FK	�I�_rS�'N&�1�a0��OI�9��Ӆ����ヺjĿP��� �G�����|��]�)"�)Ȍ�E[���]�	_J�&H�\��D[?D��TA~�[F96���}��"M$��(n�dNqx�Q�i����+qK��W��h�܃��c�Vԍ[$�A��0�z3?p�\?�Zk�v5(�0%��6���U:i����&e�#� y�Ρ��D'WF��fI�!eb�����(����++�W+�ѼQ�������D���֓���p�cx�y65l w��Rk��f�L����]���?�M��K�E `5s%Ϗ��x+���E�&���~7�}Z�E���A���Fl_^�.V��8�)�^��Gɧ����W��&J�-YcL)A��=>�=b�������λ�K���oR�c�M46c�8�+!'�N���N��r����0Q�BS&���v_kF�E�;HBIFS�a�^���n���/��4���H��	qs]h�h���o�]����d@t������_�6N���C�G\���#i��H�Ӆ��,o����ʠ�E�t���G��Ե���� Q��Ս���� �N�ۍ�˦��qm���V$?��:�:gAE��6x�
?��}�7���ړHD�t��a��)�Ay�5�ݻPlp�����.�N�)0�|�2��y�%�i(��� 'ʕ��]y<F�2y:��j��Siʇkw�ǌ��a��Mw]Q>��$E-L�A�-CK��ZN&��$e��?G~~F!r�q�^�T�-~���̎�?07�`@�O,�L;H�6���:{�	�O�F�]Q2dV>��`�:����JWM�7S��*�U�N���`�{�?dG�ąl��b8t�ʭ`�)�tvZY��&�£]�S{/����U=�y�-�j}�׽���3A*�BN~9�)?w��ـ42���"9���.�8.n��ۖ^ XI3�\$���T��LΙ��*L��()v���r \�+�II��?��<�����;�-֠����pb֚��%6� ��CV#� �~�%f���X�b�{�����[������agp���D%�']�$x������K upϦ@Cv���u���h�:(���#�y�'7�|�XOZn�T����-��A�3�t��U�6۳��#Hp�o�&��(|�@��ӆ>sů��� �^�yZmJ�����k�$� Q�zt�g�:Q���=�_�pĦH��h^Bj�쪢J S�����{eb����S�i���*����i$x��Ł�Mz��k�cL����b���U���sj8����t*���%�`�>[�QOxĎohkK��3ڡ��yD���=bv1LF1���W�O9û�n"0.	�z)�c�U�u��v�-ı�����#~�BC�֛��7q�p�KRgt����-���G<-~WG��-:�oh��e�|��u�*{M"��qI��~V�3ad�iNDH�ɞd�Q�]}@�)a0��UI:q�;��9\�!5v��� �ֽ!ܕht`�388]�%�ʶ��@\|��e������(��!�����5H������X0�ڂ�%d�g��BvKt��|w���'�7YV7&Q���o�u{�I��Қ�@�!\;�B�Wkn54���ar���L^5=�t������C�l�9_CE�O��-1�ѪK��K�ڱ�T��n�]�z3�����*�~����v���PrE��e#�2�5.}R�Mm-���}_AaZ���.Y��������Y�Ve��SD��X�qQ�#���P�ј"~�?>F���^ #r�z��9�e��I0kYb'�:�7�)�dsE�w7&Į�,kp���s2��T��ŗ��'6ş��cU~.�"��I�S�b�**SB��G�Lt$H�;]���B�
Bˉ��v�>�r������R�iMB����۷ 	ׯ�2��t�F *"�I�!ܺ<�K� �"V� |
2�$��� �w�p��%�R���CMv�����J"jE�b�ď�?G1'�B�G{�0�G��#���*K��"�?���?T��6�?�M8�UH/~��59���57��Or?k��3>O6L���D���M�D�(u�(��:��fr�K:�!��V��8��R�G�]+,��i��5�3&�0Pp���<:u�1���+ }��|~y�� �j>kx�ӛ������U0���ЊɄ��&���al\�4ݰ��CƁlY�0K�����췳U��~��
���X�s�*0K�?��0�v��/M�d8��p�9�l��cjj��;��'H��ɾR#�Bh<,n�ҙ91y���s�U"���Z����GD��r��2��c�vSW���)�ΊD��:{�}c�R��F�����?�K�+�(rb�N!��a������3:[�LӾ^Ub���2訖=Qq�s�_���ya�k�N�i�/�<�?FQ�џX�N���
i�^�co����nyGA\�+#�C��K�F�7���gl�dA���cTAl�n��~5�BzB��6�"����1���ZJ�Q�V����L/�,T��ߤ_?�-�O�
�{��c�i*�\��Prv[EB�a{�ߚ!Pۭbq~�\q���w�B%�����8�A���fh��Vט��RF��Y��H��f�;�)"0f���栢������p��2�P�$�?7���C�o`@���&�B6]�<@Kc�xfI�x?�ц}}1�9U,	�$�<�u���u:>-.�L��ᣞ��|M:��1n8ls�b�<��-��R|����x����%�Jan��
�%Ww6��}�ѕ'��9���+Y�q~�:1'7���y�CH�.�`"�\�1��&`Ȩǣ*Ӻ����9���ݨ9Z�z�Q7@$�F�x����w҃��y��#��Q-�m�u~{��A�r�P�����%R��O@uafU{x|�q�5,�wqG��2l(����{/�	W^p����0l���}�Ml���e���9�5�0���X����t��]-�#z�4z�mw�L`;"w�לY[��Y� �;ZZ:%��J3[%	�����6ƕȊs�g.ފ��R;9/]t'���6�b����k�W�)�%A�}9n̃o�?P|Bi�Ơ������V�bT�-�c��WW��*����6t��3�o��IԨ��,3	嵝v�9�Y�^�^T�5�%;��Z��:��cR+p��YC2��)"R�%0�+>d�Lڥ*N&�H���
�؋�F�o��H�j+��<��7�i�͇�Ryq��,�T5������P��nIF	�_�!T�*�(U��n_,�ۥ�F�Pn(mC� �v���w�f�m�U�1��柋a�֩`�i7Ó�w^�}��=�a�i4��N/����k����!.=O`:HS����dE���m���F�0�&�Z=^w��y�����/rZ��(�7Z�M��=��Q�!ܟ��F�#�;<����gL���d�*�"�z#�g���)��E�^��|z��^�^�b��Q^̱P.�����J�ʋ���}ܻ�8��}�8��Ti�iG.����9<���Fpli����3X?���FY�aB:�����rz���!��lq��C�*e�f����e��Z�^�Xϴx11:�"$Sz�'� n��>O�*Hd��2l���<�q�<Ú+0G1RT{�-㋶z��EW-{������/Ԯ��.���blA�q{�K���S�$Ƀ�ϫu�  و�[m�io��\���Ĵ$��9��Mւ�`�$��XzM�mu���*����P�j�Y�aeBXX��b���yx�z�%%jY.���r��c�?�#�]�����-B �%�E�՗�T�<��Jxgk�
�M�L����SU�jܾ�Z� �������"�������9��4GSB7ߜA;��9�eͨ�BW˛��W92K��O��F�<���Y���cz|��?�$���Î�ý���c�]�(��i�A���}¢/a;9?藨հK��f.׸%j���3�}�F��~�� �<K�8%�B��'�7A�>��Ԥ��;��St\0wC.W��#��K�W�E��zއ�8��REq.��A�c�	���-��L<��xJ6H��]ۮU3TML�V{ź����3��f��K�0�ĔG���'���[.lR _L `���9��\�j�I��(����ӭ4)t���$q�@�a�	� ���n&��Њ~D�V��ݼ�v��e���^�e5~ݳ�~=�#t�	A�]�=	3���Cq�ى�w��7�ʻz�xD{�	��WG���nF�)F���G�L�7��\E]�p�,wG~����WL�g���ೋh"tI���N|��k���Cn��a15�P�2߰ Lτ����)�s���¼vߤ	�f7�7��+��1Y�Z˾V��𲲔���_����E��gS��P�7�l$(�Qq�|�O����� �����j`cљ�'+LO
�0�����i�8�h�sٽZ���S������|�:˧�A	��Db��hy㮅��rݗ��aj=�?�ԙ/��+IA����'6T7 i��qO�6{-�>�R�~7)�0���0��o,1��B�������\�!���#Xb��P���?Z�m���>�r��a�D?�B��x���I[1���3V�I̱�����L�&CW����8&B pW$P�r����&l�����1�)\����ѽ#!r��)�A�i�L4f���S<�MV��>ۆ}ht�V��U��	��!��zy���kS�nt�j{廰����i��a�RD[4� �'�kh�	{��Ź�/�!ʢ�<�5^��D.���@�Q��o�r��w9,�k2�\<�=�/�vIΡ�8��9��%*�������v�o�[���w�]��s��=�a_�N�G��2 ������9��.��f��S��紦��os*�>[L/�߸#��.���� ɠwݪ�A�h�g4�( ��G��
�9���I�A=�� ���\,��޲ �PV�|��D��d�_����|B�{]ks�ԟ�݄�L'�O��4�8���G�0F��zs�1��J�5"�!����҂<�_�>O+5[ǘ���{;��-�0��-"t��VDƈ��V�8,�vT��y�Df���-��z�M���K�/��k�@_����+~�|� ��[\�M��K��#F���c����j͹��1X�q_�k<�<R���%��(�&�����6�]��<+�*e�<eok�w�;��߼�Z&�H�ؤ������nW�o��KW��ܿ�j��Ĩ���@�J�i7��	簃+J�eל+�4��2��<�,�6�PYqb�1��P���	�pkB��ư��Ⱥ	k
v![���������	��NB�ѐ�ׂ�Qx�_ y�e�?H,��[s- �+l]Fc�q���/��s��(q����"��3��Q�/[t��Js��O��o~�>;�*�#}��pn�s������`�r�1܍��~	�S�������V���dO~Ò� )g�v�<��wm�[}Qv����=�E���-(��?�Ru�Xˋs~[:)u4��K"���2C�F��\��s�~��/�����	���A4��3?����8�Kwx���YN/�kl�i4Y��^p��;ia�ϥ_ �	�jҠ�G9�S�+��$e��!��۵1�h����W�C�/�&/L�͖�ʉf���q��{J0>DO�\�!+�% M����jZe���0g�`O�41��ym�T*x�kL��^��GL�s_Ȟ�������0D���^x��xk��g��#�Ñ���}cI��YN^�o2yn�E@�"K���������MM��-Od�C�A� "d�|W}�����-�W*�Q�r�� �<��.��]���Q�3�T�]au�zu��1�?s�x��0Ϳ��Lcb2X��)�gX�U�0s ~13R4�1�s��+ZĦm�e9���,�/�}��=mN<���#l*ڼI�,+�M�ٔ�h�4��g,Ѥ�5��}�y�G�i�qO���b�,���h���]r��. Sj�s3p�p/�Н�-۾{����m��7�8^������t,�oZ�e��kYP���R&6���n��9S�"��02
L�N�����kOi�e��J�U?Ȧ)��<��(
$)]�`��1D{Y,���pN�r�&lO��� �@(Ya�S'�*��1-�����|]@����=n6�riK�Ș�ڬvi+�D�m�҇�q)��&#�jvq�M�!�CN+�)bP+eN��fR���=��c�
<Ǚ����*���Grw��7��D�ќ�ww�z�P�пy!�{ӸM����*5TwH�*��iZ�#w;k�6}~'Ih�쏀�<r@NRfD�<;;!�_����?7�j�c�7����F��yۓ��/+xT�c�o�j����kZֆ�J
�k�_q��l�v=��G��͘m8`��������c�+��f7f��V=�˭E��FT�.��k��څ0�w��,����ߦ)������['�?�RV$��C��y�E�hR��h�8�$�m$�޳��a��1d�z�E�;�9j����D��H \U��m�{���v�G�����I��H";� �H�u&#7�v;�`g�ny�?��$��}��2:M�!������-�x0��HD��*/k�2�2������߻���F�h���M��
tJ0n$�W���B��w���D2�o��ҮF��?����Գ}\�\��^�8����QQ��;!��es��;��24b��XY��9�ϟ�9U';��� 8(�O���>���!��-�+:�m;a�W���\�$������oDRRgm=7:�]� ��*+a^5�Ad���IV�	�D�Jpt,��K(mԞM�^�ɂ�����}�(g��bnL3��g.��7�
������t�y�����CaV.T A�o䒼��T�a�~��:�Dl��%�Ǵ~�w�éc����C���x'�"�]�{m��f""O�
d]#�5\
�8��5�\\�+%=�y�m�fՇ[�[d����^2�X�tzr��S�w^�c�	����d,Ee>�lb���@?�|iD���>������W�O�E�b��-�yVA����}IJ��[��mz�����u=�WWNc���󵑔<�ئ�왧�Cz�A������zgU.,v�V�D���'�#�f��	E��h!5	ހ丩���C��XB����hd4�J?�����a�;'R�%iφJ���zB��-C3�M�p�����1X�9�e!H��v1���8��q����|Ko,�4����6ػ�����e�H��m �'��17�nCA\<�ҧ�����5~^3O��s]t�].��
nn�n��}U`IL�6=C?a�ᅘNLG�E��d0d`kDl�WE?��@�@�JO#꽵�ϱb`�~�M	�Pχ&�{�x��I��V
>�;GVn/�FD	LˠV^�v�q*"�߬P��R_8#٥\wiX�:;K�9=)����z���B�C��c�C���D�P~maΧ�Uy�_� ��K��Q8�j�r�����wB�,������X>�N�]�MLZ}�< �<�P����
J�>I��B�t�&[��%3����V��Nqѽ/��y2[���K���%��H��w[�'ٮ�H'W�jh����ﾼ����SUCcP�����m�W��hׅj��_�� q/�l=\�^�[�O��9!�{V�<=}���x9�Y&���p�>ۣ[�/2Fk֢^E�Э����Ah��Y@�L�O�e�t=�;��*����~\�$��C�y����Vxfc=U 5�~�� ���E;K��^������~�|ǧB��V����&�|�N����qτ�<w�̻���oj ?[o��T��X�=�G�ظ�S4��}6t����yL*j��a�OHl��|#8}��J����a#���#�lW��TK@��	*�f_�y��`����!ˋ"�h���r��Y��-��;$L�|g�>�f�t��q��Y.��ќe��5}�%�N�� -_�h�u!^��ׂ)˭��I>Y�7<�c}��|b�$!�8�(�*U��y�d�U,t��(ܣy1�q��9`�G��r�;s�����6��f���^�,a֐��k>�s'5)�n����\�]Dޟ!!ҩ����$�|���O0=��)[2��H�g	�����<t���@�Q�"*΀S!Ԥ�3�o�.�;W�F��#T�ue>AZ3%lW}�,K��t藦=���_��881ҡ�G;~D5q� ���?�職���Dy���Sk����Ib-�K45�d՟��_31i�?�;O<"�m����6a�Ju��e ���3Q��@`ɾ�}��M^��f�/�iw/2~����%��͌3��z���>vj�H�ʜcVw�g�S	�vu���V�&*q�����?J�K��CVbS3�Z�D�a�,#N�tj� �n{m9��g��������*��E��dr��y^��L���kWt���A0�/�G������m2�~��U����6*	\���&�#�7F3PB���L7G��O���q�~z0���S��>0������.5� �<|ztA?�Y��o	Ջ.��ݯ�䟤�5�\/�����ݿ��o�!�����=��_:W���վ�*�'��躿BT��j�k�'v�����kɲH���wF��y�$b��	%��ӄϕ�m.��h�������X ��Ϣ�Urg�0��w���L�g����g�P1�ޭM))�����y���m#���)�8w��ݳ��'}#fx/Sz�{�jba�BP�a5`K�2� �ˉ�\]�oa�C?:4��dYp�{�F�A��z��� *�c��}R�3l��u����"����Og���޹�{�*-K��~��^��3T�A%����Q]�7��2#���|�1\ؑ���O�u���&MK��1C̥]/Gp��Vio����zy�6Ņ���b�!�ý=Z���Q������=��N��%��"&^��X��w,)9��uF�R�T��C>��,|ks|�$e��Fw�CC$!i����ы��1;���f�ŧ_�����^����`'�����X.;��mh���TU���f�S��)���+�ǚqٓI���6|�Mk�)tGбx^��CP�#�nTҽu���'��&��4v�v�N�v��Ad�!��ax�ad�ad������D�m���*�A�/�נz)J�'�'��sf"��$�m���a@@<Jd�I���݋���^�P�}�ܳ�?�����/:m�;w	�m	;?��!���=Z�2JT�k�L_��K��;j��St�Y������mtL�fz�h��8I��N����OM����2�M�)��"���'���vH9�d�y+�7	��c_�G6q���.���3���fa$�7�Q�M�-���SZ��Ew�����jO�x�$Nb=(���?��,����ZΩ�'˂O"<�Y5�*cC(��mf�:�f�z9�Eve��L�W%����_�M&�6�U�fX�E��ms���k�[^�z(���u3��.��~��.�ɨ�!��������r�M+,V��7����O�#���o�CQo�z&4D��?y�t���b7\	���c��;�ja]c�T% !9
�eG*���`#o���W�{/��f�4�lm�*��-��������2D���*��]��y �g�a��R�b��Oc�|�_&�^K������ �KF$�iF}�јA�����Un#��u�"�&��ήV��'�O#a��'I��k��
�ۼR�c(E}�9�[n�~��m��ӺL5�,��+� P,�M���`����H�R�07>�8��x��Ѹ�� ��,̗B��oo�M|���j eiK𡹃���	�_u���[�u�>م}���I�[6��n��|��A�R��*2~�����?l����s��O��!��>�o�+uh�"�(�@S�Q�ͅ��ᓺ�K�1�#���������QB�$�J�����W��o�7�����no6���{����}���{�5h����d��4k�x�u����Hh��Px�id,(�i��?�i;)��9��A\v)����,7\*���S���<����)�9�����zv����[�5¸�ƮgɕG1�([��)W�^�"D1�%<�&����_��|B�Tu-���zBx���������T,8���V���C���,�8|w�TdL�D�5"�$��Z�*�B�z�&���.�w�Y��9#O(Aq�'�qf�e]�;���W�]:�	��?��#��_b��1Sʨ�Js�"�N��b����
aW����t��tw���r�'2��3_���=�ye�M�&����Q,C
=kyR�]|�u���ݢ�j�����<B�ǡ����lVua������5Y;<�EPC��πn��A��?��.nk��P_�a*�!��R?����
���0\cŷ��Y�5/lj�j�;�P�@���/���Z��&d����pꮟ����?}~KT��C�_}�w��lƝ�gV�J�h�{��r��نP1��p�Gq���/�V#%`$�`��겔���ߴ��*�ɻF�d�󳍍���u�2082��?\�"-S/�j�չ�+�t�ޥo�4\������j�w���
O�������
d,"�D*���3�2Ǟh���P�c��H��hڦ�ӈ�����!���v/�v�B߳r�(_��!�'���N��!����҂����i]V���ݛ��؈��Ki��>!�� ����J`��F��n�7�@��R]N�6]��a`1���BV"�T���U7���(QϽ\�e+� ��ِ�ֲ#��~�C�?���?�[�=���a��%")��1(qz�.��x	1zny�?o��}V+��K\M>k�h+V�I����pwW御�4���Ӣ�;1�
R�F�.X�vj����8�Y����㓄�b����������F�0��<�'��_+�Nw��K�oh�i�]~���;;��P;Y�n(^�9V�h��(�g���n^��~\��T}����7��wд�k�m�(��E\g��y��ܴvU�WI����/�<�<W����/�	��ӣ�����T�Ry8g0�G�'4ӟ���PQ�"~�+�OUz��hsC��� AU�/u�ڸu����F�*��������gO���o��C֜8|�*���T#~,(*�2u麇���8I�	0ή�*܈~]���dxg�(�TV��Gl���� ���u��fJ����@h������M���*Ù\<��A'�T����$/]Y�`�]*4��['�j�2:�>�z��ujp_����tf�gJ�p�3�������o�$��r4�ɨ a)���R���k�U���4�wު>��"n��-�~	V��S�5�{9�m�S��~n�����(����ȠqaIl�i!x�A|��>��Rpk'�� ��b��y�KI�Ͱ;�^�ji�g�9��}C�1?�IS����+�60@�ʖ:�(����rx1zӾ!�^(�w��ΧԸ��b��S@�pr����)�t�� K������3�Ԭz;o�OI'�{�3���妍�
�ӓ8CK��3�u>cʔ�s7:W��.ۯ4g)���%b�N6k��K��{N�������d~E��{��Ln:=%d��8[1=
K�ME����;	�_�Ǹh�ե��OP���'��A���ꦲ���4И��ث�O�>�a��0y_�d���0�e��9���!��}!�ST�/f�RU ��X�'�ͧ{J��/AG*�~�ŕ��!̲ٴ�L��V.,�N����`���� ���P���X��x�N�A�M�J���'��i_��}%��C���D��{Q���d��K��/Z���%؟�M��yex��5���.a��߲�~��$��6
������.��KS�G^��W�?�K�>�~���=��ۑ��a,�r����~2{���	_X�0�P��NA����	�1��8�O�g�4�_p�zJ��Ǔ�������Ԭ\��i?�bZ��S���K\E��U�n�L�擈�����x��=�H�M��\m�~���@~`��Õ�g�i�_�"�V�L�����r��m�����=)v�����H�q;Ӭ	�~
>�=A��57Τ����:�'o�1HU�-< Z%��z���%۾�Й�- BX�QY�їP/�K%�gj���O �I�`���g9�` R�x��A��"�L��{�	M��0��Tx����s΄=.Q�T+�f��P������F��w��ĶRZ��n>
Ǜ�G$<%�
��U?J����bT����(�isM��o��~��}���*��4L&� ��)f��#$/�]�H�s�}1���ӓ��y�9�x��6y�_5{D��'c�!�;�mb����nɖ����`��M���rM�]L�����<(Ȁ��1���������~����K�b��M��V��)���L�ȔDI�xG,+��8��>�N��4:���^I�Zo�G���T�Q\[p�5Ӟ|��>�����<)H�1h�?��t�P���^�V�)>>38�/�<���WV�z��"�V���ͫ�E�*y�xʀ3`?\��r�	?�#���ؘ�|�&�ql�0_��ȳ�)�͐3�=��\=�����f������'�5r�8�p*e��&���WM&3���n4�ƥ��=��EU]���:���i�3�Iy� �Z��7F�gH�	؏+��2�̾cbl�e?�%�hu�6���rA���6�5��."ؠ�/n�\���ٳ����y���ޏ~�e��m�f8^�����%W�uTI�
�2��|��d�W�7���Q#�B����W�vӉ����9��--�)�։ w�٦ݥ|�����&��S��*
�<r��4���,ɣ�+`J�7�	L�"��>�^�����r>ǵ.[�X���Ѝ�D��XJ��k4�Mo���˓��C�G��� ���վs���>맜��Ǎ��x�ݞ�gyx�G�<�;�k�>$fؗ���-�	>��G�������c��Qн��x�hx�n���z�[���祵?}4st"Gi^ƿ����>�Ęn�!<*�i���ѱ4�D����G]�EIJ�7�-���k�`��^�U�K#�t�
J�4J� (�݈ HHI(")��]C�
�%�3�0���=#���_n}����ٱ�Z�X�\/lY(��7�O�|�FZA.;�w��$��e�QwV�"�� ڑ����F'hL��u�TWU�{�s�+��qG-����t�g/AަJ�	�T|O��g:���Ay�,)�(�����ܿ���
HF୽��_E��p���R�j���O_R�OT���g��>���1g���ݜ�9�\�I�� �e�������-P5�!����s���R1�c{&�r2:M*�������2��h�����C~�?��&Z7��E�m��)��>>	OoU7���Fg��*U�/|���yn?	r���G ���c���/�Xј��zU�Ϭ�2��a]Ef��F^@��W��is�W��Miz�s+��lB�.����cSF�z%=n���CR�An�����[��nug����]X��F��dy�F3|����1�.B���1j�������nW�%Ⱦ�iZ�9�y��>�^_A���[������דe��V]H��X�t|��ZE��Kq�dp������iⅦ�,�)�!S�U��@�5��8�F�CT�m�r��,���,��?�b�gb�ˎ�.)D݃�l�_O�Y	��%WO�1�\��BD������f֊�Ņ�/�e���Ҵf +��O�4����k~�:D����Cʫ����W)�\*EU��\��D�j�&|�]���KMy�͔��m�{�1*��˗�e$��;]�qmU�alg3Uݱ��,~A��5�vp�����Q�e+_#�pc,�/Z5������5J}[M�<��y��x�OF��\6U(�:����E.�')VV{�K������M�S ��iva���!�o"G��@��YF��O\o��������nq!���P̐ʕ.��\4+ox-��(B�~;��˄�}` \U[����k�TEI��y��ˀ|������77�#pdJ'�Dͤx���K��ROFCYdFy��!c�I����\�PI�:A,bqٌ�ht]eM�'ϭq]I��٩\�q�Gj;\�՞��Jѻ�=?�"��+�����v�"���~yC���U G��=dK��.2�����1B��~D��{�U���'����,#!3�Ճ*�����rt�\Ԇ`ݻ� Zm#�@R�
�0[�_�?��J�.��Qj��e����A�:9(��db��]�u�<�-}iyp����&6�?b��YM�: +��G���wD/b�r�Ju�s~sͷ
�'�2oq���L�5��e��L}��F���8d������q?����.�#�����6�������Mu۹���_�>�f;��h} '5�y�*��*����������H��_������n��
����lw�w��7��	3��6��i}��k�2O�3e�u���N�����:����"m�vI ��Nu�7����w�s�L���)��C�V�PB��[^yr)˗X��zO�&Ȍ,��U,����p�z=��չ��NÞp�rd�i`-S9����^Ď���r�aVS�!s5��4�����,~����i��wK�eR`� ]���\��ت�^y�L�E�õ������ �z=-�z\��aP��iH�� �\�U�1���ׂ������S��S&��531��ĕ9���ޟ������z"�2���Mv���U��G���Ow�~U�Bۑ���4K��D�/|�hj�]������g���a�����/���a�}{�O[OI��g-��s{T���g�nʴ�y�Z��^�&:��ͱ�Q���+c���[z=!mw�𛿱1�-����T���&+�,"F�t�3���Z2odo4�j��F��ӄ�XxD�����p��͂�i�Wp��W��� �F6^)����c��w���	��$@��}�1(3��7Yf@m��trr��ڲO�+�/��ZrOW��H�r��?][��j��+;�q�y����g�E/saG����/��_L}�Q�Cit��c���S��T�����`!�4ѽ��}�l-���u�Y�pB���]8=��>|��a��ͥ����}��gH��1A�W��A,vֆGG ��<˞��l��6���т.�+��yջ���w�[� h�/�U����⫧sn�N�M�ʛ6R�ͻ93���߮H��z��_̿�2Jس]��`��s<d�sW��3������9Y��ֹ�M9�����L�ҋ�x��� �C���γ��]�����I���9��R���j�@ʗ�Fgǃ�J
33}��s�z
�����k��8�z?g777L�455O�p�3���"��I��)E���k��F���F�L !�`��@/�L��WUUV8�z���8�C�����#� ������$�Ȅ�@Y8�7�k�$��dS��p��[ �}���L��:�U@���%�� \�OL���Y-E�����\�ę�,��:�� H����7jr}�@�]��ۇ��>��!���&��f?]3.@+m�n-3�,���-�4\�[���B���&U�Lc`��"A��h'��JS�SE=�y��'A�:�T�?������~������s�X���>����Ʈg[�E48�Z��`���ÍWq��H��W�����`���x��V˕J�}�N�9�Mo�	��%Gx��)�ռ��(��3+`O��Ҫ���]M�Ϣ~��Z}�y�<&p5������/fT�0��ߣ�|��99�z\N����X�X�u�I�gx��2���_����z���]��8��<<c�*_��5���թ�`,�� ��~B��Y i+��[�b����@������}!�S�0=��h��D�)�0���׎��A�3|��SԵE~�<��_K<^�D^��`�����C��
���$;�fϚµ����}ĽN���K�.��g�$���6��V���q���s���t0�W��Q��g^�4�&��a���r���3��i��ڴ|�1��x"�64^X���m��ϐ&>`�j�=��x����jLC�WCz��Q�D�v1�-���ũ�kG���wvvN�:� � CZ ���fE�X��|#�3��X<�k[=�����k�ͧ_�D\�����?O��x8/�JN��0�N~�;�ڝ��[��ɣ��Eq��)-������8f��<@p�| H\QQ�@J`����@�l@�>	-o�� 1�i�H{��4�X�;��UYt��x퇀Q�K�9(6��������q�����;H�L��*�Xz��LMna!WsK��yFX�<6?L���E�����2I��T�!�@�y`d
T��:ո��kl��p)dɥ��M{/��f��[Vѓ��Ǆ�����jhX틭��~���y�~�+�T_,5/>V
3p�Ó�����rw3�z���m~Y"k��֝gg?��{A�k���wW'QF��!���W�+ͻ��Nm���ߺ'Ҍ~��)#Ԅ�52��~0��R����Ih{��X������x:�ڲt媤$�:�����PB�x+��KN��
Rͫl�.V2�GL���|´�9w�YA�m��@ʭ�D�����a�?\�[�2���?o$�5��l�>�)0n3��h?���:��.��o�(m��hw�)��P�G	@��~��^f/K&��8oc�b��=��V6F^� A��^���1 
@�[�/�uD��|���G&���g��K==����� oaa`�oS���8�Rt��?HO����3s�Jmߤ�`a&`ΐ159���mx����lfB�fMol���f�L�3��:�����:##��j��L3�O�3��TJ��G q��1eg�6��(�����t�K)���{8&Wmm�_/@�;D
��J{9��dq���ބ�[������v����?a�8n�qo+u�M��T�Bn�y ��o������un.Մ�5..�S-�jF=$止[|ǔKݻ�7:�i�5�@����Mc������������7H�O+�*��Y��ζn��:;O4�&�$�P弘PŢ�H^e5y.��(����g��s�,O�&m�pn�5�,.���s�3n���J�%[��R�2���kz~�شl�8��Ē��h֦�v��Cֺ���~�Z���KRc���N��Q�0�u�������v�U��^H�e-n�	�oxJ���^sm��rrTd����M�g���6Y�W��!��5c�����H:
8�q�b̈�3�1�<i�_�mEf[�-n�O����ɹ��f��� غ���y�
�A�*�����Z���H8�R�҆4`�3�v+!�8�M�|9���,�"P�W�Ld�ᒕk�\�10hZ21�r�X�)��/rq
|����h˰ޯ�´B�m/�����"�)���.�KY�;���G,#�N��V}wd�
����~ʂȝW�_�FX��G9ۿ{�I�RGD�Q�A���X_�r�$�̥ԫlJY����|�r|p�Q?�hU��u��C�i\򳑫��*�L�!?h�U\�O���m,,sm��q���J��E����ҾK��Its�#����lW/��1�8�������?P�y���M�2]-��s�nӬ7���>�̽W�gNa�/O9���m]ʠ����������%ޤ��z�;� �ޅ��Y��v�+�G�I[
<�b19(ʴ�nwC�m�R�c�'C�;D#���3J��B�cY|��o�ʋS��f��ϛ������3y-�OieE>��L$�юz~�{aO�*h^���-�r8�+K��0g\g�|A ��/�� ��K7�� � �>���mh�b���� ����x.��E#�k�>CR��t0ا��Sʮ�`F'q�-��?El��R[�>��]�*��΍~�d�[�	C��x"B>���,�����6��H
GI�5���O��}*~���<�q���#�[�,9q�r�K�nd|������@�����K]?l%���R�Z�*'�*�^f=�����5���)Y^����?�\k��߷��T9��q���P�:O߂��d���"9s��?)Z�~B�Uvϟ�N�6��	�&��2�w���v�r�/��*�9�X#�&r=Th.l��8D�,]�d���y6X�֢�Gu��T�ȁ�H� ��ʯ�p�"���)�Y�^�j�^�.j���st��o�	De���S�������4�mVr�.�B4������N.�=�Uu�ߛ�����k�`�6��? ��uD�P�j���B�em��.�T�3b�ghIRjv��n00�
��wH#��i��s �Q�j?k��%�V�(�����#Qtm��ǝE�W-�4��JETĎ�ϼ���Vg�Y1ί_G@����Yml#^9e�3oT�c�
2�Ł,�����J;9�3�hE�] 9wO�~���f�*s�b������<�W�����ͦ���~��

�d5V�E�iv�hme%�	fP�"pe�|��gqŶu�E���>��Q]E�$����Gn��BaV��� ��R�6���ry"b�%�yl �P�t�-/sD�:;۽"7�ZX����Yj�k1�����4*�T"M��P�wZ� K�b�\�j]��!aΈ�ð�Ŕ�*��a?������~<<_rdPN���K+d��"X���Om��-��?9���ӹǛ%(We��9;Q/����DR^�Ŗo�*�i}5�U����|��H��o~�P>��5r��j���X�`�gzX�X����{?�����#���w�J���h������z�c��}�n�{\s�B�t&�Cs:����j�3�'i���)dA�o|�0����GDaM�'�>R���l�M��̉�[^�j��8#M:9�T�����P�Dٝ�>����#����{�!0?�bv:z���(��3p���X�kR��E��ww0w���G0ݠ���z?c�|냜q1�h 4�66T���#Ng�A��l	�u�ϒ���>��`䂆/'�%����t�k�����3�=�ޅd�=��4׸>���6kP��
��}�y�n�g�g���0w�0�{�}�I
�����XX[J��J|i�c�=�SI�O�ђD����^��k$`o%i���'�<�(*-_W��K��� y��aE�������9�?'[��NF�$�A�J��*eB� K��x%�>�y���msP|:yǁ��૥��f)1��>�~�c�i�^�ت&���	ϫg�Az)�v-�@��T�Ydz���<C� IFW�[��䠵R�%���\����i��߭I�/7a��PH|����]���g;J��T6�t�O�n'��"��/E����>�Xճ%'r�i|7�|��_Y4���PT�%nc��
���S>,�C챩bM�L������@Õ}�eM�/�i>��%�$ �3}�#��o�m$5�����<9��9ڱΞ���S��M��^��]����*,%i��vs ���~g,  9�����f�b�b	{�٫�"�E,b����[�R� :U�ٺ�疯o�9�H�����N�S!�T�w�����W���>&����w|��Sd��Ծ8��Mc��l-
��
� �%2�WY�ygb�T#*�0��l�{8�G`��H̑���3$����
`��2�<���z*�+� 䂓 P��ް/?��btJ2�	������.�"�ڀ�bҬ(��4�m��F��d3�Cy?�j�NF�f��O��Q-ЛZ�}B�#��L���޼
�5�i#n}�҆�:�CښPh���ȣ�L�|\��:��(�Jv�[Z���g��v��)c:xiy�,>��<6�W�P�$Gp�B�(Uu���/�ǧ�XOe׸�af�O��6������k.
��}
Ծa�\=�pL*�����=1W:������$D�ʣ/lxr��nk�����'�yhs/O
]�[��ޭȤ�E�Pw��i�}�/�1��_�0��0�U>{��@V�8�l:�s��M��?<���H��B'w��&3��HĢ�w:�m2�t��u����L�Ibn��3[�gKy�����:9H�%@� �Mo�/9�s�L-Q��ܙ�T�J�=J���8�}�}��T�����'_H�Iu�RB�����}>4� ���D+pG'�2�	��yR� hQ�������x�g�I��#؈j�` o�����y�4�,w��������Uin��� �1{����"��/��%�@f��|�_�N�҃�;��g��|�G>�8>���C,�����7����\�S�	��Qi^v�[�ۯ|��lu��,��n'N��T����f��f���_�SaIĢG��ʖܑ�I��#�������SG��^�]r?��|��}�{�
]�����s�z��%(��/Z�ο�mݴl�JӮ��y,BZM�|�����k�����O~Y�}�ĥ|���E���ј"->�Ҧ�m��)l���,���?7#b����]��'�h}�~���{AqmNB�x�_bҤ*O��?�Lp����NV�}_�{�(����r��dȜ��џU$�gvg�nڏq�Ѿ�퓲���xji��u���	qYA ��3���X�����;��^Q��>� 	:h��Y�Q���Q3��b���Ё��NI�rIx;�EX��g���+�0v��~���}���,�5CL�;���?[ �Ҧ�m9�>��8�A핞�7N�oR����z� FXK\f4[���l��u5��3�T2n�c1�!������įDwE��Y6�"!h��-<q����#9��{�j��Z���$t����!��օճv_*}Y����'M��X�L��WS�����
kB�A1�7H����9:6�bW�<�o"h��CN6_�y�=ZH�k"��vG��R��v8�]W\;z�Z�U��ǩ��7��&Χ�'J�$��\�\z2Z����6�+���L��G���6��f��C�DY��R�?{��,r
�`K��a,�V��b"�S	?��+�-�+k�� [3ȸ���������,[���u�7rЗ�8|V�����{���r�o����W��Y͜���X2�����%�uG&i)ԙ���B���R	>�|��4e�T]�B4w�q 9��lX
KL��G���
_���e�r�8'tU�Hye�o�ZDWz��h��v ֑x����	��>�i�X�@#��&�J�+K���r���a�<#����J Z��Z��JX�k�*�}�&������dnr`��;K�52���ƺ):���˛|��.LuJ��u�Uz#�M��=�cڹR���L�Tx-�O�~���|#; KA�"?��
��^L���3��L�f`�]dy�L{�M
6��v$��H`��BE�f������H.T��L��ݚ��c�奨Xp����.1ќ-�l#�	DX[�_�w%�K��"��|s20�~I�(m��v���������h�����^!#2�*Y�V� #�3���H������c<~���	��Ġep�)/DKRr����Y
k �=+J�J�t���[�h.wH{������	ͮ�e!����-�U�L��Ż�ݞ kP�eޚ��fYe��.�"���O��XFv�����L7�A�lC\����H�����-��O��+Me�� ����rN�g�¤��N�;��$o�˚`�R�Tʎ\��:�����iO�}�w��+Ow\�T^�D8r��֬�9�_�u��Ӵ��p� ����ך�]�Ybs�H��s��U����~���lg,q�ʣeZ�%}��W�1a[+Z�A���Z����)���f��iQ�R˻��v��'*���r,ؤo�5�Z������k;"M��X��e�U0K1�>��|HNĬ�3�^G�3��[�5��1��ŉOP��e�}���7��5~X�lI�3�Y����X��$ʡ��]s��la��`���W�d�0���&"w�Mv�wI��p;a��+��1�����97�s�iu'!�Y ����.ñS��������fQ��	+H(�O:�?�Ӱ���B{���]. 9?�y�!L�l��jK�pɗ%�P@���������6���KU6�s�?���,��9+]qi�]v7��Z6H�|��ǔZEz�S��jI������t�cRrԚ���|Ź�X��܀�h������*d+��Z��ʾ�(F`T���69�j��t\�A�!�E��T�[���'-T��\D�t���-/�&@9�̴`�^��V+���R�� �����Q���ƖP�?��b0��əb��;E����#
��Q9�G�e���O�K!-W�)�6L��%����������|+w�N����Jg�A�R	k}�}�hۃ!1
��b�,����O�sdE-O	Z9��h`�����Y��3b N:t�{����"&��j�78�[9~�_�o]� iG}��#�(�k�Y.^�%6��)��o�����fM��_����'����6����
�7�� ی)���"��K@�CSS3+�`ϕ;y�����k8��~կ�-��ꝊŅX��u&�˃�e�6�~�*`|�B�΋'���,�g���z"�v�X�$�O,�m���
s���pڏM�W7��ar�Aؠ������U�"����p5�bz�.�����"��r%XݮEK��-s��Ӯ�g���C?&�D��V�|!c����b�UP����I���f|h�孵1�����y񋸫�;��fM8��O�5�7Q&<�O��$%�;�z=Q�ez�p
���Q:.� ��:U;+	�Km=)D��9^�Q$����۹�Kr�8�	k�S��t��5�md�&�z��A��;�5�(TҳP$	�`#�6�J�n$�y�R�4|
�j���e$�8p����TQ�淌�?��D4��fw�޽TKV��|&�O�&9n߂eXO����$Uw��Pi_�T(�Ҿx�葖N8�[�}r�,����q����x�y��hA6���dЍ�_ћ�%WXe�'�����5��c��P��f�A�#RAR�L
�&
��#�(8x��Kم�J� 
��tk���(Op/W�11�j�g1���9�y�����Ac`�G���k8Z������ɂ�g
/��F�Y�������X0B6E�*ƣ��l�#�A��N�oY;W�cNn<Q��_m<%s�f7*z�T�3*��b8�SQ�o�A����.+SZJ���$�{�]i"�ͺ� �Xw�C�gF4Y��L�R�B�?��Pз��ի�Q�����"9x�.���;�����Eę�R�;���xM�v���@^�Z%Eg���\@"�scij����A�����]n�\�R˃�HE�,֙�;��Wޞ�sA�t�<�{��t�vh�[`]cu�����0$��w2p���_r"���~�3��@�A�8(��T N��-�7�v�>o��=�ZD�9@����H��?�r�J�p��c��b��Ə����������m�V�@�%:saz/�?��v��,�e����=O��ҾY�E�8�2������:��ވ�1����e;�<�&�]��k�g�j6k��o�Ȼ=Z��[�����ԫ(A1&�6Yv��_~���q��(q	����zl�/m�.b�'C��Ǯs�h��R���h.����+2��ߏ�<N�姈u6;����(Yc����)�dY������X�$��??��� �c%����Y$K�·Q�����0�y�}�y֞����l����+.8�G��حd3̎�aa{Xق�Qk����H��v���&��!�lK�h�7?ή������������ſC�G�܁�2I��H��h�pC 7��+��u�a�6xX��x2�m'Z���WC�O�H�V6�����z��@�)���������<�i ��9t�"c�zO|��-oVE΃v&^�|{�c������f7؜
����?8�տ|�o�
ؽ+c+61��l���{Q��$�l��Z�g�,B Y+=�X�N�a�>�x�TZ#w�2*�@����b�S�o'"V�{>S�������Q�ءZ!�9@w����x�*'�}�aMV}Y���8]6!���ŗ/��X����`�������]%��K�1�T�E 2r+���]Β�a�Є�x�]?�8*Dȥ�cw��
�J���X*�k�� �OE�wr`[�a���FE�Wx�g���5��FX(&Mw�r�&���t�
�?B�4��o8/���e�@�d�|��'���Rf� ����
JT��X�L.#6[���=���=�_�ìv�R���}IX�� 
)G`:0��/+a����\鷈�R���y��D�@Q�81�n�_N�cp�g{,d�Zᩐ�>Q�+	���C�;f��~�-#ώ?xN���} _�˱R�~`��:�7��bFg�v�B��
f��'Cᑦk1�k>�!�v|x�l(�T'���Q�L����N�����*��d�xq��ɿ+����U�1F�\��m~�P�=�ڗ�?��w+ "�ޓ�����R��"�j*K�[@���#�^afgXΛ�Lb��h^ܰf��� r����R�&"_��a����)��JGk�&��d��g��u�I����@�r|nRa�@e Wu",�k�������$O^�ڮ���Û�u�Y&&Y��I@���b;���c�R�h��y��>�~�P��2��v[�Td����ѷ2#�M�*
���P�����UϗY�kʛ�k��8��u�{m�~$g�r��T`g�ѭI.�@��_��'�Iz̼#$�@:�5J���/)i�Q�e�.�司{�s��<:��XN�� -�߬����$o���M����mN����~S���'�&H�{$����pG���x.a�DI�F SbN��{uy�C#�Ng��dJ����3ɂ^�.JݰEv,,�b�<}NTjֿ[a_`�%,���&�3�:�����*�Y���@�_�i�ݺ�&sN#�1"����kq����H�&�mA��Z;�vU?���}�>(K�ڻ,M6i�����iKߐw��e�,`��i�|���1�F051} 7�g z�?O{E�����M��]������r���͘ҹ�~�9�H(l��2q��8��|��������@�t�g"S�dm���Gз�r�w�z�X��*�q�v�/�#��%Ȼ���L�Q�v�>֧������ t��c,.�gA�}Ȏx�ލ�uJ�{�W��U��a��/��W���$td:?��#��:e��1f�r��ؑ#�u[�GK����v�*�d�Ĕ)I�B�>W|p�/2:.W�{�u��2��8�H���v���:��-H��B��������I����x�(!�
:LA��z�>��<�e���&�s��������� �l�a�'nM�ܬj�W�5�	�	@B�Bz~��;��C#�8�J��YD[�*�W$���������0\�ή�m�#
Qd'���P��t�[K��_)�N�%�1��O�PZ��� HsEQ�#��'|ҳ�t�����u�@����t�[[�F�M��;�(�:y����Ԃh�S��KS��������Lj��[s�+/ ��"����5"� �n��\4�?_���hԑ��2�+�WMW��wW��;�yk�aRz�y�%W�t}�F�n4?�PT'�a��k�*�E����j�'�O�I�!1��@�xeQ~�Y���&FR�P�ϓ�cC���]�')������������!�5���c�5\���y(�k{��;$�NCl��u����#�Жp��dA��0>m���#�ۿ�D(����R�	l�bIZ�Y�?��h��l�מ��N�F�S�w�!P��sgλ���I�������
z��P����������B���[��$�*��RfOo�$vO4s�d�{��[�L���}R>�X�����{!��k�{�#��4�Y���Y���/���eVs�"��⣧�P�u�bs[��͇��j��Gn���#��DC��y���!�y�aH����hJ�L�r�h�1u��,r8K�UD���!�)�w��X����l��B>��1�u+A��D����N�$���Φ�3���bSt�x�p)�z:G�;7_�䋫�i�}�J��=�WV��ڣa��5!�Q�7R�Y���JX���S���Vux��-B�n�L)�.?'lՐ����XQo��ЩRߙ��p�/`���3܂)lPp��	4����q�S��L�
�/�T���O�.��P��Gʂ���
(�]�ϹO_*f����F)���Johԯ����xb��n!w`A�N�R�XlX��F|��5u��:X@��E*���0E�U�$�T[��>o�ԝC�	���_�� fN��r:=�ƎrWГ�(*:�V�~�ϱ�Z�T5�T�
��~q&I���ؿ�a�M�ޚ	 �(�������?�+k�B��<���jG9z���]�'4�:�e�$�ⶱ+FwT������$�-d*#��D�X�R)!��C��rC��I/h ��;*�f�ۨἙ@��Zfr-˶zFH�H������S�P�4�}�xc��[@��:fg�zU�-�爏��P�&}崼3N]���y&ҭӷ�i�?F],_0��Q]�o�؍�/5x!b�u���S�ς���׎fOE$.�?��~�]�ӑ�߯[/�S>-I |l�����_j���pͲ� ��4���#�T��3.�9�9_��@�/�i��{x2:�5���p���c z���Ѕ�l{^7,4���z�v��J�in*y�A�ǈl��d����֕�}i���㍆ϐU�
*{��z��`iK9
�m�o�Z�ą�fs�W����E��������x����S
�yһSV[)S:�M� =$����<���L���Z�r���dg��b(�U����ڞ��٭ܝ_yo+��b|(�ܛ�QUfu�������JN�`�gqFm���Jzv�7��n}���K-4X�Z��6c>0+64���Ҍ~Y!��s�tb�	�L���#�y7�(wD�y�8���sYLy��+�J+r�.2io�
��-\n�h�i����T����M���*��+Q�Að�WP�V��&�si؋6�3�AbrTRbFlGE˫�-�s*<�z�)g;L��Mv\؛�ARP"�	�{�,?��v�>�ɶ
g����y�;$G9�r�����D�'\��ә�Uz��L!����r?Z��;,Cs�.�q�Q���ۊs���
?~���A�}]�F�y\)����L�٭�����B@?�^����w�t$L�Iu#�����������0�������
Je���8�8��$�N`���D��Ū�å��K.�w/�T{��K/�S��&^�\_��圿:M�8��ԩ
.�j5c<���7��,���ދs�ro��7��3<���]�' ������dCb�&}�R�۩`�?�HKP��x�A*"��HS��Ty_��o��8xw1/�p9��M&}\Lj����{
�m�Q�l��,��A�C�\��ᗈ/�Q��	��<������T���e�Y���6N�d`<��u˼�i�~�����b�l��2l8�����PTb���քxk0���LSsarS���Y|Bk�W�a>��F�|w��� 1���qS������߭ZG��G�F-U0�V��Ń�l���ùX��K�Ҵ��Eq%V:���jߧ����+>�@���{���IϤ;N�_��G?��x��ԟm�NJf��I<�� 5˯�e�~���������>�;�?��I�q�����H�"J_�Ł��vގ��ſ~�r���X"����w�0������ºe^�A9Uݲ�a�w9�Q�K�br~jD�~�Q����v\��d�˪���t�F}��+�c��\�|)�Ŷ���f����|�����Q8�TO"���I|�p�<��G����H�E
:&���&��?�^U8�O�z^�9>�>M��Nv�u�e�=K��(SH���5d�p:6_�v i�O^���X,A�baIj�b�g�?���ө�<'t��L�H/K��(��' :E����7v%�+��ܘunPYr�~6kq�ᢿIݷb��{vj�>�6���Xllw�A��� �m쎠��GM_'��?�_?���{]g_������+	�u���0����	$�zSiA�	��X�`�sYX+�ǯs�Ϥ~ w��a^��<�I�%�p��7��Yi#MS��$k��ޗ��5���?�����n;a2�111qc���#9s(���;;��%f]jW ���ܥ����e�|����>�f��]�S�Į���N8>*�����y��4��>2�I3�Q~O)P+.�P����%
�E?����ӵ�"� ߗ�,��g~N�uq,D�?'�m�Tnl3Y5G'��o].�j����w�b.G�fҖ�����çm@���P������ӡ��{N@��[eMM�Bڎ^�,��3����]���·e*|�s^#e^�m(e����"���"]T_wz�4[�L�܁���߈+D�<#���x�H9�4��:���$|����ݳ�Ҹ�<��o3O��K�E�ۍ1[f��g��Z�&oTnϸ<�T��cU���N�W�x���J���8V
'בQb<nV7c��lfKLm��{Ă��F��V���'�͞��W�O�oI�Rԓn�$��5���ӞFY�>��	��y2��d5c����b=��s�]E��e���������byY屮a�4���6P��%ft =�){b *�_��:{�⭣]����U�C^�͇��$=r�Ҋ�8ïKvCr���{�c�>oɔX���n�U]�ý;+�m@J�5k,D�N>uylJM�O�칹a��,omÑm�����Ny��J��K����y���`�`�.�埽\D�+t1��A�Et���rp%?��l��Eb��/�n���tT2�-���`5�^A��S)'��V�"�)�;�h,�İ/��6N �7.�,!��,n���GF�)�&��>��W��t����';�A~�}��o�Q�ƽ��3����D0�W.�ADBr� Q��r��aQßƳA�J_���`D�Bۙ��ჲ ?ηo��%�3'�?	%%G9��q���=�Hăf�#Tߺ068b�[I��n�#��	�\�D'.�9X$��cݸG�p�����(:vsʞ���y!�*m,:���z�=�A�V�f�FR(i�q��o�t�6������,����PU�֗�ϐ@A<~~�S=&`9?��_���^Qn"p���h-RD͑A�����Y��c�4�kק���oA��;��E��f|q�0�i�!���6����?�h�I�Kе����[���6��X�6���%g�r�Pv��j�^B���C����@�R��B[+N����3�n��J� �:�%��ӭ���oor������B�c�Rs���0N�V*� k��^�za��v����D�t�>��	�9N�,`���K� �&�$���5G��hH�#���'K��2�����@��3+P�p���y�e����(v,��o�_���¾���r+��/��X1W�#j��j�>��k�-Q��)��1�N�y�aA_���:�m�>���׭(b�B�E�ܰs�9����W���n�=���n�V�lg��!��yeq0�����hrZs���_b��ba-�guJ�wF�Pq��W�r`Ǫ�FB�(��������<��g���� ���dU$����c������u��;��u��JR��M�w�fCA�]�2�B:hӼ��V���g�N��2C!�S6��R��rz�݇�6/��L��s^�
T:�t��q�TC�/����4�8�ɷ�#	�{ycY�L�ܴʵ���B�o%=�x����y�a�_�gVz�	{��Jq�&��76%Au��Γe�f��*y��+J����ޛ�C�v��/�R��"k�v$!�v�J��mT��'�蝢��(E��}�d�:�Pc�f�f,�;�K����������������s�s��s�s��^���_���J�����I��ƴ�:z�U����7�����q���!m0D��ݮ�蒖��c�m+����-��7+��1�+u[/R"���7?J��9����������r�L7YU���iV3��(9
{���eK4	ӑ;�j[�@���gÖ��}����Ӛ�E�]j����Ұ���<�-<��w�p'�$���	���cac#c���x)ϣv5+�O]jf�X4N;0�8���29�۲���ڰᤥ�y�,%�S7<��M�xX6��s�1ګ|������I��שּ������W�����ː�&��r�]#^FIjGc���s
����uι��׿�Ե���Xf�����s�d4wE��g����U���1�����~�~�yc�9�W���skKNn���2c�pu%�c1�N�HA��s?o��c��3�*�m�z�ޕd�3�,��#�n���>��[��[��b8?z��3�ĉ\w������_l�.f<O�g���B�/|���M��۩���췍������ٺD�ܗ!	�{j� �ӫ6�Q�NML�9�_�Wr�*�f�is�I�����]��D�U[qf2h7��c�"���@��J:>yCx�`����9�/����.�w��pS`�>�G����`b�C'6�W���;�^�E�Z-VY̭�w��JF	=���9��\�`�]���'��5έZ�~A�����_�T�|��o���˿�[9��f��+�T.�M�y�^���%�mj:�����cOC=*�<4hǚ3���b�K������������ ��g�W?�ѬΝZZ��(�)����"�o�-K�W_G���b�鷞�O-�>%��n_O.��y��.�ѝ5}=+u�y^�/s;�d���˸ysv�Ȝ�7G�G�W���S/�d
b�����oR|��Zj�m��9���+��:|�Q:-7����_H�-lq��~]�ċ�W�_y$e�L�ڜ�Q\�Fx�=J}z�zۅ��� c��Su'
5����7_�q/������>/�� �
�L~�O��V|/��I�umEՎq�1Z���|;kM/Znuk_ؘ��R���Tt��|���<a/LF=g�����0ۻw^�1��>���mҾMR;�ʙ���q�C��Y�22�a�̤ꋓ2����Եl�]U�X���=Mʜ�EnSq-%�Ѷ���%�_�yP��~p�h-�zF���
�Lb��N��	|�n��^�l×xb_�I��;���خGR��_;��m�2կ�%,f�i���{����ޭ��n�������օ6��cY��2L&J��!�}���i<8T�M�΋<ZDiu�$�Jo�k�)`�._����ܥ;l�n�OK[��)�O7��X�g�����D�c%
��Ԕ�{
Wg���UZ�՞�zc���W#{�9�ch�������?��s��L�֙z����C�����<�ff��u~������|�$Ffc �hڴ/�u����P�z�&֟�m(���)��9ɛ�ǧ�Ǉ�J7*S�+ޅ݋�h�­��g���Ͻ�e{�BOY:^�%�D�4Pƽ��N��}�1_��r޴�X����E���*�u�D���&_,�w%s2F�G�:�:�ޏ�V�H�+髟�[5��>|e���dw�Aj��)�8�[�|�O����~�����,+~�7Q$���/0�
Ͷvb0Z�F��cV�ݯ������ӭ�~��Ԉ?�on��B}��i�d\�r�s�q�}�E%�i����4��Gj����W]���[Bw�����b����D8�a!��5�v��w�V�#��hˀ���}:.Ǘ���Ɔ^U���4�J�}˽�.��)�y\�@�\����p�(F�1ổό�ֿ�e>V>0����4��묤�y��d������O�υ�=
�>q���zR�5��nP��zV��۝h7���S	�}�KD�)�ǧN��#.\4DT������;�m���|[�@�O��f�ǋ
�{S������?�A��xr�u�I���~��Ĩ8�����p�۾�z��и�b�X��l-|�}T�Jyf�\�(��[�"v�R�vD>�~I�H���x�k�<�$�PT�kB{\M���B�]�N{�9]5oiRR���YY?�a>^#���QL^�N�'M[�E]���:�:�g�����6^oZ�r�y�'b��aY��s�.�X4�,}���ihbK��w��y+��n|�>ʵe#�ofO���&�a��ΰ{��>h �L�>�>	E�w���n�9���6{�
�o�3�x�L.��wv����7GDb�]�z�a��n�h��3-���΄x���.�/�ʳ��jVa[X�.�<�,&�q�	����M�s�{���s�aq��a���}Q�O*6	��n`���T�d��5 ���WeW�
�	�<��{�����ۻ���g��Q�y��p�������[��[��7�3�G�_��Q�*��;�P��_���z�s��g�C��E)Z�Q�o8�J��eS~�Z1��o�Ck��n�NML�ۅ��v��]�d�_y;��6�SnI�A��7J��K�Cj��1��sԖ�|.��Yb�y5�"߃��__�ל������O��Ӊ�R�#�E��Ϋ�ʧ�������i�ī��e܎7�b��Mc�h�����myg�6�7��hR�D�,l�^�����S�l"��j�_�ϳ+����&xwj�g�v����ô?am(�`��	�]�񦀐�}������ߺ݇
]�M�����ɠ�h���g��O�8��+�?s�z�ݪ��9�ߪE\��w)��9c�7�0��ϟP	�O_�i��ƣK$o'^xh�S���P�zN֮�|o��.̒ߥxw��y�\�%d�i�H��/و��G����g�6?6�b�.SYO'����wj����+r���=�<�홱�K�-�Q�O���s8Ɍ����Q�cKʳ`�Nx$�g����������U��#c6�������ʡ[����v�K{L��)��Mt=���܆����$���ك0Ҫ�����j�ɟ\�;+s�b�SG/
�,��mU���V`Wf�������>_�x���iv�.���_{�V��Hm�K>����j�qS�����+冋�4t��t+�Ժed:�w��hy!g�'l��JÎ��.v|���wb�/N��11�q֊����=�Q�6��o�vM������ҷ{������&q��^q�iDA�8a^��>�������և�*W���I�T��k袘��Ч�,l������Rڷ9����i�&����wO�ND}r�{>g�9z�i���b��D|Xe��J�7�=:��/jlx��!y�x���r���=�7�YR����/(�������������\��ϧ'�vPW�����=ee�t�x����i�~�-&��&��(��/�p������ZZ���9���a؋�k�Ԣ��͙뿽��4/��h,��\������'���VR�Q{/��Z�IJ��Ms��;.��^�)ǋ�>���c����g��]5�ʯ��L�c�U�>�j��iv<P)��_;QW�n�?�պ��n���%G�I׾���r�iK i�����}/VR���C%�:s/����x��1g	������ôiK�h�/�����oJ����)�X�9:u�{u-v��pF�s�{Ea�7Ocٚ�9>��M������]y�8a0��#L�hʱ�o����NOQ'o��.�����S�z&P�~�2]���l}��F>��,��:��S�W�7�U���u�V�@{!l������_6C�+z��<�V�UⰧVR���h��ܫJ�B��ˏ4�q���|0�m�aȾ�ݦY�Ǆ��)��~sNȸk�(s�Yu���+���z,�]���|8m5K{�H��Z+j<C��9���n���{<M�X��>���Ǭ�W?)in��]���&�w�'G�e��äx���;�rb���!;�,�{=l����}�@�\�IW7�}��㇬�����F�����SҿL?�n�5uַG���uu]mZb��.M�9��T�zj�f'9�^4����B���P�/��x�����I���n�@ �Ǒ N�2�3iM�]}��l�UM�*q�Bڇ��ENF�:�{��o[�-m�j�j�~D��l�fzJ ��鋧~�+Z"���wv����w��j�7�#� :�~�a�Ah��i����D�+n^��Cw�Y֩�����u���xmh��[�D�o_�ft��H����J��P�X�D���!�~;����Ry��{����M���ڔ����'��G<�Y%�?nlZsm�Z�'�\�j���{�Тڏg��Ҏ���W�?nM��ˇ���yn��6U�vEF�B����^���T��?*�>ǣ�&Ls��D��ģ��'��`j2���g�j-N��u�z�\^l��+�0Jk�����n���k&���7����T>/����k�e�m,k��*�a\�^�w�~��yo�%�Fn�K��{��e�<N�%��O�V4��n?�\e�d����P�=��6i�>��,ǔ���#���~>��{�ޕS�#�G�G�)sJiM�m�վ�����ΩՁ�Z7�Y]i|?��v���}oXaY�9y��O���u�7�m%"9�G�����<��ϧ�N+��t�MN,ʌ������_��#n<��l��N1�l�ٱ=p��*OK.�8I�y�$U#��N�<�ױf�i��*��oy\�5M�s	�~<]�){\�t�S�C5�uO�U����㭀���C�yJ���������A�+�ۄ��=,�_�r8e�v����q��Z��o�y��V���r$wqװ�j�q�'��,�\T�I��\X�l�|Fv���ւ�L��.���z�Zb�r�Q
ơ�g�m��nX���9�r����m�����+�]
U�t��xS!�v���y�g5/*��ٟI��yɹ�|܇zi,+�'V��q�}�e�Pv��f,����,��`�Sj�m����;>7�~c���MYⷹM��~�(��z�������s����S��j{P`e�ʛ��)G���0��=\I����"~3�n<b݌�3�L�tL�*	��T��������z��\]W�<�(�����^�������?�:���xH�P�u�T�V�*�oK6��T`#u���̭�:�m���h�]9�X�aE:/q��F�grL-��4яK����'X~�����䕯�+$j�~�<PV`S�z�巀߀�E��N�\�a�g{&I�_�ϻWǗxui�L��g��Jq0S����l�!*+<9D�UK#�B:pz�����}�v�ҿ�<�:�3�c����"��e��p������_Yx���XK߮�����g��iK�?����Z1<��[uQz����Α�ŏ�kK��iO/W���ݷhI��v��gf+7�T�d@��	�~��4oQp�e����E�n��Gm�U�X��Y������d=m���✞�V"�QV���νg]@X���Uz��Zr�)[��)�ȁ�h�f�C��.-�m߼8Y�k΃K_%�ww�"�'�~�p�d��C"�b��зCw����*��/b���w�Y6�����V�S�g�X�0�حԾ�*w�����W��H<U�#��wa�;C�`����s9�F_C��za�����n�O�}�p�V.�Ӕ(�T�YwC�?1�E��oV���9��+Q��48LZ0q�	��֓�U���#�G]w����*�׾G&X"���󔉏Q�0h�Y��S8�A:����TT�ٷ��<x���C�o�o=�}��C5�SQ��9P��=	��*_�<;r���˸�����j�+àw>��+�vh�?V��Sn�>���<�\0��9����u��EI��}=^�=�cѣ��︝y�?٢|��`���w%lҤ��N�����,�A
۵$n�݌��94�-qx�S5�p�BՂ�\��&���W�`�Ȗ�m\���zk�M��O����}�D���o���Q\wZ#�];'��8��p������V0�z��{U�Ò���
F<Vڻ��m�݋_*'2߯#�1WB	�%_䵙��׾DX��>vŻ%w����q.�J�Ej<6@��y㺮*˛~���^�#�x��-凛�{�3Ft�ɒ]�^.�崙V�e�IR:Ń�Ld�:<�j�ߦ��r�U7�!�պ�J�asS�q��7��?�xb���Dq������o?����݂�'ory��܊�6r�I�%k4ɍ�D�x�MA~��������_a��d���ݝ9��5�򫬞��c�����t��^�Ԏy۵�ڪ�:���H�Մzm����5]r�C�X����|]X����;<��>+������ɟ�*����Z��Y@kJP?2x����Y��2�����,J:�� �:��?�t`*-��Ӕl]�azG�`[��K�&M���t��X����O��͡��ބ��=J��_rM���FUKb�N-���?�T�`?YW���)p1Xb�?c�ܟ3,���g������W�NW�j�M��'�.^f*(�w^�?���XU���k~�)�o-�ǎ��1,O��1�ʛ"�b���c2�Q:[r�{�h��_�"+�}Mјؘq&Mc��-�a�kQ��N�[���bsE*��o'������|֦�=Uje��S��8�����his����֕�W*J�
�jj�z�~��d�%t�6���EG7`�<���&�.��bYLx2g�{ұ]�:��/������7)P~25�Y��u�����I�������;�gH�z4���"~�s���?�jv>��#��G���n4m�xt��������\�+ϥ�9O�~�kH��>��ٴ���O�5��怟Ϲ�Jκ�C��E�(o��mO�p�b����V�<q����?�����F�%��.�U{6�-j��{�r�M��VEo��{���-k�)ɿ<����[>s��T����x}x��B�BE��&����oW����\-���l�C�j�{�0�],{Q�&���%\�Z	�d�Hϕ6�n'�難�MJ��!R�/ރj\ZgI���.�s����s�m#+�O��7~�i9��c���h�/�d�E�CԆ�^D���N��i�ɋ��8�~��7����\W���7�\��b<�Xy��
N�v����מ3�A�u>�Z�ɣ
�����)0��,=h/ꜻ㜤�ܛ��~��-���:H�a���1�[L9��;����pFzK�c�=���J~S'��q��b\�M>Ƿi_i��&��^���R��� �*��yi��F��Ãu��i#6�Y�����l�=�frTQ��;�\�!x�/`��'�؉;?�o����F2��W�f���d}߅�;���&u�|J��RL��'�|���N�k�kT�H��5V�B��o���{b���k�+� ]Wqo._q�<�ڻ��Zb�O^72��S�-B�^h��3aRV�|u����ʊAOxP��S�4y��b�L�"�l����e��#�w�f�O��xq����hJ���I��}�o���]�� 	�D?���s�;�OZ<L�~�W����+�A�ІҪ���v\[���=��4�Kw�i\>Ns�o��yi�k.@ӺO��0�F��=�t�E���Bs��q��OMmi:Z/�ۥ��g��k��S�_L4�|�L^��k<�"��r0�͡����$�P����H�.��&����x����J��-YS�}�m�5.U�K�	Y2�D���K���/�W<�������o��
��{gB|�$I<�?Ё�S�3��[����Q�ɱ<����]�k!�1s�c׮)�u��x|&���&�u�V��s3�&6��L�5�q���#�f�ՉG;"�]�w�T���M�q٘�>�w�H��k���]wr����CVO�>~>����.��K{�2��X�����N�>��n{Ɔ����r�Ǹ{z�a�4:���*	���)��&��&��Ð������h���Ӌ����R����oL��?����1-WC��rW`�O�Fs-��7׾�<�H����r���8�|N6��vO[ p
(䍄�K�pD�*��;�n���\������3�vefO��n*�����蚉$�49v�t�d�c���Ѻ����[��������<xpN7�X�/V���[(C#T��ڏ�n���L��е��Ѱ�\!�R�B瘽v�l�&�����w�Z1���Jo����菻����%��_�'E��S��	����[��(�*�V��5g�IP���y��&/��W��)�n;���e�o����m�"5_$T_K�?�k��wd�½w�^��;v�����.<Z��Y����M�+��l&q��K?a{7�kR��:����Y��1�I�B��W�_�헒W����Lm;3�>f��n���wK}���KJl���Y���)[��OM���s�2����ύ9%p�����s1�s�0+WVVn��e#V��8�K�Ju�Q�}뽂�jw.[,��>�l�΋!�:&����ȏ��fq�CAwf5?�$��شcC�≟��޶`o'�:��6�����P��/���h,&�Z �5��K�h���xʌ�]�񂥼��o��<{*���JF�A���鈸3R��0���0F9��fDzi����T��1mo�,E�*�B����b�^Y�n��D����{�`�8��'��cq�R�)9!�ܴ��/���T,�����Qj����q�z��1J:���ȋ�M��Kz�J��MZF�b����J-5�?�M�3#E�1��<������SW���ˬ��W�Ͻ:\5�9�����k�W�t���f���kxTv}Kh
���1��������1�|sB�U��I	�ʋ[�4e��܍����ȍ������,��ӵ�J����X��0 �Pvq��阃���ƈ["zx���s��n�\�y�']u���P��I�q��;����L�(����ٙNK�C;צ�S���\*�x��ZX�����R����������$N�+���M9�k=���x�'�w3Ft
���Y�Z�ex���:�E��F3o7Dϵ�0�Aܥ�����I�z��_?��1ʞ����.�+��.⣅.�)�N�n+#.n�k�,�@㾯�όj��PFTdh��0������e���u�bo�3ք���u�1b�GtX�i��e!ACؠkP��H8k���� 
y}xb]����`���,��fj4���=u ~�#
�O���X^�P�d�F�.8_�{u�Y�������~��t��"�#SA��IvF����X�kӛ�����v�e���<�j�ؖ�(���1�4?�����Ώ}L�"�-��M�<�zW@67'n�}c»����)=��*iکup�x�:')�)�I��3Η�J�	���a���%*-#�5|u����K���
�,�.�Fë���;�0킮o5n�c������|d���=˓t�!��?��|4=��d5T�n�ƺ��V���5oL�FFds��fh,t�Do�_`�;Kk~�2zk��,�s���H���&o���u�Ē���Z��0'4|^�)H#%-܊wBesٳgy; � CA{���i�&�[�b��@�'��s���כ��|��=���ҏ�<e� V�ЧI���;���ٟ���t�3��$��J����l��n��j�0+��^ʈQ�>�2t+��$�J�#��CW��s_�� ��D!_����=J��Ҁܺ�+4�Fޙ��@�J0$ѫI_�)8�X[#���Ǩ��}1 }��d�p#�h�ff��s�}��I�*$��e�c�SO%7m�����l01N2A������涊m�sb�aa�D$����ey�?�4yH���N���?{�0�rDo��I0�m�vo�Լ�*���(���g��Q�#��W���܇�z�]�4��M��
�@|]��1�O�����ِ�جB�;0��L����HK�8k4�a6dh�� ��Ak�� |������ȳF�T�'�����Sv�����ќ�h*��]��Dl�m X��/	����k�1�ȁ�Fx���#�ťqi��q8C�hߧƤ\��^}*|q��D!#�?߇r�ء�ɇ�Ih5�۫��uS���т�U����az�BQ5T��S�6��o&!���?��x���>�9彣�Y]@>:��1iD*��Ԇ*;B� ^��E@o����s��t@+���=Ϫy�c�V�mձ
�a�ֆ���lH&nw�sr"GtΜ�����0�fD�q���X��vd@AJ�s���Bt��S�mD��[��*}O����e^����~d�� ��@|"bEY)��Wֻ����YnS*����|`1e���|r��z�6R���lj�W���8�Z��~���������X�s�<�{��:�p'����Ǆ|9�5�8�(�R��hG��?�^>�n�K@��{���G��� ~�T��+��)`�"Gr.�aj{�Ėd�i?}YiF4��:�}�ⶣ��!�[�f�}o�P(j�[oޜl��P(�P�3z�=�`ɢ	r2�]3��s�#Q1����\wv'JR��l{� f�Y	���b��/��O���wļ��j-�߳�l���٪3�@h�V��!�#橭V�>�Ě�}����=��6�Iy��ȉLZT�b�w�	A�ڣ��Î�x�IpP{,.�(����v&�=|8�-����X��J5=�퉡��6�n>�����5�ak��ຄFF��ng�=�����Mǭ�'��O%��)`��ec��|V��#�'I�b/�x��񷿞�'���D�"L��{{�'����lD�3����S�<vsߍ*�j��ԓu���(��ܩz��+U�C�?��P����폸u��G�޳]�JBv��H=8.����}�����S�A��9l>�D�<�w\-�t�#K���������"#��S\G��Z���=�u�d�r~lpI�����G�aO{��ͽ O���B	c���@��o�a�d�#��j��3f����}tƿ>vcVaVaVaVaVaVaVaVaVaVaVaVaVaVaVaV��z�?
����/V��V�.ۯ"1�A���^�;, ��w��k���:�ή���:�ή���:�ή���:�ή���:�ή�+Zw6D��(��t�|��~�vv�]g��uv�]g��uv�]�/\n���׻ �_�2�ή���:�ή���:�ή��6g^����\P�g�gbE�3驖I�Yh�&��-iJ�W�������*�MƼFtc�=v?�u��k����_���j}�bh����z�Mm|����l�g��+��mg��50k`����Y�f��50k`����Y��_P&ߘ��d���7���|K�<��-���(/'��v7���2:������wb�wI���|/����r�yc�
s0ڈ����	O�w:�������ʊɦ|^orDor���?���B���RxE|�]�,9�:1y���C�)F��0�ɸ��?��/��,��9o�FM��:i����i���~T��b�\#�{OﱱŒ%�e��'*����0�'>\ՈY)G=��-�H�X���I�*�������3T�W�| _��WQ�ĤFA��x�~�DRY����NL����jIc�b�Z؇�T���Pu�z�&����X��HN�b��е̠"dF�,*��r	>�� T�w���pib9��nvb��ɸ�_Ȱ2�����&����߅?oUC�,E�0����y��|�퉊
�󏼃%��Ɵ>��iQ�rE_��(h�ہ}����)�7���|P�F���`&Lp�rl6t�P;'I(���=�`�E%��~�O�����{)�X�](_�F��f���N�r��\��kޝ;1y'׼���2J�؜��ڠF�ܪ���&�a�np1�/ӡ�1"�
�n���'�Q��Ȱ�,M��l���Tx�(�����%��>���?�SL�u�eQ=g,�∽���qΑ��Q.��!���TB����.��$����'S��R@ċ�	�G�$� e�B��(���Xi��sl��w�nF HB��y3ԑY6�}9��t�O����g��%N�* Ჷ�s��n��#��+�3�#_~���>�3 F�#n�Cʼ��<�����]�[�!�`�𶙡0����%`�O�y�ϟ�d(#�5�9|r�)�3S�?��Kt�Iq���nHQ�*��ݽ	�������8TN37�D�!t�7����l���q��p��~Ri�yG9��Cԝ�I��2'�*(�Q������F�, "r��Vt^)�/���-�����QVe�ڂ���D��%ePbMr�T�2�&
/���$�d�Ex5�����L5z�ո�����Y���Ah���f(��iAI�1�t��oj�ā����/�d��#da�'Ya9C���`)�K'�Ā�5�#�QR�/��30
���L��ڸ��tP ��Ӝ�IBT(��)(���q��t\���ÖL�I����� D?�J5�K'�.�U>1�d��Qo\�+(�DdREPܷ�<Ce��U����� e�T�V� �ԮAҍ֙��.�+C�T���Du�#���w��2��əR�t�֔���݊	zc"lT�:�����b2Ȭ�����>��C��6�s��U �Np3�u�L���Qg')�ŏs����nO�Q ,�`41�H�5� "�5�Te�L���	FʕO'&?ч�>�\+} ���F�L-��"����F�́�-�ٱA�]��WPg�D�VC������98�﬎�B�Q����3G�w�,)Q;<4�ϟ��������IK�0lx�>s�l���������N��V&��57���!��&(7��L��upX�ߐ��d����q� ��>SC�zh��w�ߊ�0�3�^�A㜭35i��12��*]?�,7�����wa�S� q�Iy�3A�v^E�P�2m�;ᝉ3ѐ�
L��͠�z�D1p�DA_Tğ�NVf�Pј��)���qj?�r+���(Cqa?�\�.=�u�M8Ȕ����	���<�F?�PCE��qxp�L+�Mx���H�S*d$�q��������d�<.�a������o\
�#�`ɝ���qѡt����X3tdt�#�6@GF�؄7�#>�
N��J��������ѱ	�0i�DV��Б�R�<�����	�+�^�A;�� :��������ꭔ�V���̡k��Z�2����׆f�<8�C�����:�Q��@����q���KG�A�Aߔ=�L�+��S
�����F��[��鈎�@��}))�a������l�����«7�5���u�'�53t����Eo��a��T*}�����I�����|Vv;x�`�8������h�S�+g~P��4t�I-U��wH#g��ۣTj];Q��\D�}x9�H0��; mF[d���[r��	� �g� �� �_��'����n��4���.�1���H#_[Qa�1��G�Ժ���]zR!�E���O��U����Ol�~�K%B� �Q�����2�5h��-e	[�bOQ�����|�O��>�Z�'BI)·r8n�ՙe��4�_6T��Q���&�9�}����� ��^8&o�N3�������'P����g\���`hC%�}��%P�i3���@Q�l�5�m@ABܘ�����م�l�ɏT��Yd�@����cXLPv�#��CVW�2����d�eP��N�����f��pP�gtȍ�ƕ�����������"��YܸG?��ɹ��?C�S!��wg����J�C��-�h�5�!��yS*���U���ȡ�D����C>�T&���^- �&�V�7���'Ɠ����H	���ߐ�^�E>5¬5�v|�BD	Qb$n������/�|�Ռ��F�r�u'����\���F�y���7/����F�\�An�z����qo|*���$���+�9���������36;�ȫ���p�re_���:~R��D_������v�Ers*g�s����G�f��L�N�HS�D���wKQ�%�@���Ar`���ޕ��Gy�����r.�.B%��3ݐ��?�a?@�o�HmӝI%�t��oVָG��S��:@u���%�� �����$�c&MG����Q������g�~�x��b��"u����
 �9�34�T�r	�����3I߹&��1��b{��w�@��T�u�f��c��ȑ WVQ��19�}���)���:�|~/��;�zO,p�#����b$��޻�=`���zo�z������`��*��,���\4�^9�Q�G��Y�ȋ��1ȡ7�c�ģ�NTQ��,�s'�5h�(TU/�@(��J�	0灛{�I'~��M0|&+y�����>�N���O� ��0��Kj~W��$a�'�L�K;QY.���Uǰt�O �*��~ �W���Z��_3�F��@�x� Jsа8���%�Tu A�Y���p�ͽ�d�!���2Q6�}��d!��O�42@X"��M턽J ��d���s_S�׊��A(�(.�*�^&C6CR,�2l	#MG(]�@2_$�F�ޢA�Yr�0���.i� 4<��R�W�$�E�!+]ڎD_A�;�u��Y��h;��N2��:��]����J��!K����-c���"�!��%%�ˬ�;�ډ�o�{õG3$;2(�U�b?��$F�#�E*]r��fGجQ������߲�BBpݡ�f�:K�&� slD}3W�N�z+~�D~H����K��sI	��^���.)��ώNm�{��=��܈z����F!�A+�Cw*���fT^�p�3�	z%~|�	y���M�#ݸ�tIl+��c�� s����(�q����-�� �����qX'p�n�鉁��>�I؋d�H���2�e3���Jګ{=X-�[zs��Q���Y{AF�A�*�1��L؋���n{�,��{�\��ڤR/s=�HF2M$�YiSK6��#���{7�#{����"�˼{Af����D����Z���)G�"^����\�'��?��"������b��(�%��rȗA	!�B���U��2�f������-FSR3�w��@0#u&��9��߼�$6z��KfX
��RtĎu�&"�:��f�����tC��9�̇�v�._���X	-Qף;@�r'w�є�:Rż�Ԥ��"�	|9V(ƕ�(@��^��IG�a����8���蠨��h�$�1m!����=�����A,�B"D��Y,�l��� �1��/!�_���5��)���|��Y(ʖ����I�e������)�/q���;m���QO2�iY^�EV���r醌�`�����dt�T4���yg?�_��9�~��~k۝Qhs�P��Y�12Y�2w����b�e�a81;�)R�@syM�q0����G"� t�����5�B�`��cq�d3:j/�ƚj?B>4�e��C(��HbO�RC�E$��˭�' v��-*4,��"�hX�Pǰ�)u!��Fj�j;r��5h��f�Є�(C;Cmr���iY~oL0h�\I�����a=8}M�VDZ��Nk;�p�7�S���BC��Z������s�[�B�nPAִ��Kj�3=/���N��9��(�Ks �	���0I,�-u�Hڔ"��8@j������1@�����~b�0��Ajw�!���?>�f� ;��\N�I��H��U&��&�r���ć�*b�~�Xp���A8P����zp� ^,��	�p»Cd��^��l�����^���_��K��[�����(�}/�H#��؉~œ���!�~^*�sA��S��,h��\W"��,-��q�A}��Wd�w7��a3�ڋ׼$W��ari���� �]�"]��L���D��כX{H)��:N�"�.�T�;,sp
�&�#}j��R�Mkp���a/��Z�S�	8�pk�AMw
HW�2G�i8ő�5@J��"�ӹ�S@*����zrZ��7t�HqeM�c�^й(����C��q-CK�h��ʐ��A�l
~[��&4�cI��V�HQ2��6��؂�]d�w�.�V�܏��7�2ut�?��&n�e0���2�g|�B2%\c�[-#�B�3���yK���c���{�'��)�Ռ>؋dx�wܪ������\�^�7�} z�^3<��2�g~�B2�P�!e& W�h���$;���>f�}z�p=�!B�W`/��ؚa�2�fx�^Hw�M�w��e��^8Z*O�L�5��=��C�$��8��[K�z����G��K���83c_�l,A� �%���6���"��4���1hkt�}�YZ*�*��V�F,��%\Y�}�PH.idN&ƪj��&Q���Z>���A���~[ɕEe���s�K�, �����$�md�Ҙ�AÑ��Mn�NɅ�N�#�c��M��c������O����K"�2n�\ko2�[@�����������<#�!	�w��&A���B��&h�� ������jЂ�W��(m���DH!���@�f��3\�fn�� ��e˸�P'�=^� �N�8IL'�j{�n���B�A(�^�s��'!��pԗx���9u���{F��qV��X�c_���I�J��C,p����]�2��B%�b%Jˉ��:�-�F��������z���<Y繲Rz���	���1(R�~��bh�3zWAoٍ~0\���bYxy�37G@�&�b�߁�*
��r���pG�.�sWֳ�����y?��k�O�E��`?�w���rsą���%�2D�I�X
QO���|�C}���M5s*ʅ˭u0�|-�:�0R���ڶ:!�C}%I�R��\��-�6�ؑ^�+��g�Ok3K���:�D�#�B3��Ϲw�Y���y� �t���[��[qcB$��>f��������^�'ޮOQ_��<Q�80�E�o��Zd�+�<�́1�Hx®#�����a	0�+��a>ai-��E�p���a^�e��~^�m��0{ �2R���f��L�$���90!�Wq�4�V�K*��i�8�S���B�r��0�?�������p��'s:��ӾB�T%吡VѨ�-Λ�SH���:$��>�"�
�>������,�H"p�2��V�3��(R�/�G,����A2�~�xH�w����J�*��'���~��$����%��`j�^����
IR��]���� Yx�O`8d0�,��Ӛ���u��Fh8����\�k���[���Dϣ��W����-�㋨[�}�+Ε=_���D&Ae�!��	�P<!�'!<<�����܈��U{�m%����֒�� d8�_����|(��3�6E��[�Z;�3�Ǡ��!�>g8�{�nPc�!��N�A�((E)�f��j�sGw��!T�<<H�Kkĉ^uB��7�-u� ��Kg}QvE��f���X|�s�(�-<���_ο�w��";(�Γ:���҂���M��e~�/�
��{������J�Q���:g�l�5h-P��xi輦~��F��f���,��#^����rYZ^��يF�<nP�+;N�E�\��"���@��A��=UÀ�[e��F�z�3�B�mB 4�`@�g�A�N|C�*���ĩ8��,-s��-�K��{��b���rnD4%�4��@0��|�^��ږ(��
-nY�,�3q��XZ�H��e~ځ��f!W�g-#�>
�p=5�{E���-�ӎ�e�Ұ��~��g\O��'9� �����_-|/t�F���[8�p�p��,������O�$�U�����ވ��0x8�F�t���ކ��^gY���kv��/�!��B�����Ӗ�v�[H��Ar�vnD�h�!E���E�#B�=K+E��y����zrT����<�^g�ۜ��M� �G�F#���FYێ����Hb!}Ή]ڡ��tfs�3��K����D�Q��J�ڐ��(,�@JG_9�r��"r6j������@�1�"� ����#ކA�)�PGצٲ�e$���XQ��+��b�E��r[�sO��9��>�=�yϹ�f�n��R���:f���g�A8�3����Ƨw���s#$3B�N�_���Ƭҹ+�O�W���@<��� �2�* &�u���UR�w˅��Ư��B��)"�I?%��g��{͊��y�sʂy�CB׬�OȲv�ID��c�aD�����R�O\Ԥb���W�6�����S�^���g�z�=���E�B�7�j���a^�R���0p���M�WlQV��*�K�?o�>��{��^�g�
Y�Z?����9g��Ա ����-ɏLH1��A�WZ]n�M�8�=�]��0h��Xh\��
��3|D@n�o���u)�jd�i�������R�O�!��t����Ъc!j���'�-�x�ʜ?z�ڏ�46;��|<�������p��;tE��p���t���f�_����nu̖���+��u�ަ�cs����z���9���T�0�V����<g;b��V[Ƹ|Y��6�a��QY�$��x Qev-m4�h�,�@�q����S7!5��g-�7�h���̸���dÌ�cxo���`��|�]K�R����º��g�
l��3<�+�Sf2+bhU�Q�4�zݤ��+�_��u��Z���R�a\1H�����"RC��~	�R����ٰ\������^O�&$+n� �Ld�b\�,\ i��)5�J_����ŤtJM����f����P�{�\o�R2t#�e��ܪӆ��\y�a��];9��g�PK   �p1Y��g�  �      jsons/user_defined.json�[o�6����k������ɺ`KV�i�n
�����J��"�%����Bw������(�����C�����I�il�!�yQ�,�&ٺ)��]�38C�L�I�[���χݟK}�>{Ye�b�nrM&g�7s��7zmo����?9/׶.�zR哫���m��i�t�d]o�4)\+�&'��X�+@� 5� B�*�8>t��6�.V뾷��o
���(��c�
@1N�&� �9��\9[����Te��i�\ �5��J�]/�)�I�S���׷��ʽl��F�;뮮��̫��!)7��E�Z�/�j�1Aj�$!��v�����]s��=��MY|ڸ�*ϳźvcؾ]{C�m��b��`�+4u�Y�(�����j��n��:���/a�u:G��pA��\/�G�ח�A<���3��~���Z�[92�� A:���;��t�3�.z:d�t�s�.��aBD��A��誧sM/I����4zM.~	╏G=G�ɱ%�|��^�G��K�ku�UTE�̳�0�-�T˹�^=oW� �n븘��)�x?B4�3��;�\0��^��̈�TL�kQɻip:��}���O`<?���`���燓�5�Z*D���G$���w�B��ix��5,������0�5,[,bns�0���"V� ?B,��0� �Dy8���Q@�CF� ����#�p _Ĉt�LI|�x�{8��b�˘��Ut5``+�uQ��G���n�)Y`��Ni7]}���E���Ww��V�^��q���~U��\_�j��o��X���O����H0��ei��b�7xU[��ڬ�1@�c���l϶���aHe�Bΰ ��b`�匧L���=�:�a�aP�#�e�4����B�୅3)l�C|���ףP��W�m��}X�~�<�U3���y?�iF�x�WO�Ù�O�<a8�oU~�<�w����>�Q�I��Ćf�[|�P�S��c�6\��9{����c��/#�v,;����W���y��X�Gʂ��Ύ�*;j��^��8ƫ����1�Ne��׈K�){|��F��K��c���1eO��֨��Ż�Ǌkt�x�?Z\�ҏ(<v`�>��i�J�~U��a�r��{��+����Ⱥ.��[�]���r�
�}����.�"]����~�t����}�PL]nrm֛�֏����wV"1K������O*��K�[ǖ�l[�g�_å�dQ��EU4�{N�l��{�5!(O� eҀT)r��Jq��w*���L��"8Ů^�ݏ:���a)%:�^S�z�lW���q�uΊ�)v&w��t�bWpc�=�5�Sv���X��>�۲�3ُ���8!���#
7gw��A�`j&0�O��!�?q�<:.@7�?.�-�.]�#�׉�M�cn;R8� �,��H�P+���03�s�{�p��9�y���?PK   �p1Y��O�K  ��             ��    cirkitFile.jsonPK   �p1Y8�w���  ��  /           ��x  images/0392a38f-5b07-422b-a303-6a624800f9c8.pngPK   �p1Y�N��i/  d/  /           ����  images/3825b8ca-e3cf-45cf-b79a-668c63877d2d.pngPK   �p1Y�?HU!  B#  /           ��z images/585092fd-6de4-462f-8499-92296fb2c536.pngPK   �p1Y(-�� 3S /           ��3 images/a48cfa0d-8c50-4ef1-a8da-0cf94db079c2.pngPK   �p1Y�7}b  ]  /           ��>F images/cccccfac-78ec-4b9a-a64e-108b6f3d2b7b.pngPK   �p1YXs�銙 � /           ���^ images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngPK   �p1Y��g�  �              ���� jsons/user_defined.jsonPK      �  ��   